

`include "uvm_macros.svh"
package wb_uart_tests_pkg;
	import uvm_pkg::*;
	import wb_uart_env_pkg::*;
	
	`include "wb_uart_test_base.svh"
	
endpackage

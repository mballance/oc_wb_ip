//***************************************************************************
//*                 wb_dma_infact_4par_sw_seq.svh
//*
//* Copyright 2011 Mentor Graphics Corporation. All Rights Reserved
//***************************************************************************/

`ifndef  INCLUDED_wb_dma_infact_4par_sw_seq_SVH
`define INCLUDED_wb_dma_infact_4par_sw_seq_SVH

//<imports,gen>
import uvm_pkg::*;
import inFactSv::*;
`include "uvm_macros.svh"
`include "wb_dma_infact_4par_sw_seq_scheduler.svh"

// Class items
`include "wb_dma_infact_4par_sw_seq_items.svh"



// Forward declaration of callback closure classes
`include "wb_dma_infact_4par_sw_seq_callback_closures.svh"

/** Graph Parameters
 * 
 * Usage:
 * 
 * Pass parameters to the scheduler constructor in the body() task:
 * m_scheduler = new(get_full_name());
 *
 */

//</imports>

//<include,gen>

//</include>

//<base_class,gen>
typedef wb_dma_multixfer_sw_seq wb_dma_infact_4par_sw_seq_base_t;
//</base_class>

//<graph_cb,gen>
typedef class wb_dma_infact_4par_sw_seq_cb;
//</graph_cb>


//TODO: Specialize the sequence with REQ/RSP types
class wb_dma_infact_4par_sw_seq extends wb_dma_infact_4par_sw_seq_base_t;

    
	// Test-component class type used for registration.
    typedef wb_dma_infact_4par_sw_seq wb_dma_infact_4par_sw_seq_t;

    // Register this sequence with the UVM factory
    `uvm_object_utils(wb_dma_infact_4par_sw_seq)
    
    //***********************************************************************
    //* Class Data
    //***********************************************************************
    
    // inFact scheduler for this sequence
	wb_dma_infact_4par_sw_seq_scheduler                  m_scheduler;
    
//<item_fields,gen>
	// OFF=0, LOW=1, MEDIUM=2, HIGH=3
	int                                              m_gt_opt = 0;
	TestEngine										 m_te;
	wb_dma_infact_4par_sw_seq_cb                         m_teCallback;     
    wb_dma_descriptor m_t1;
    wb_dma_descriptor m_t2;
    wb_dma_descriptor m_t3;
    wb_dma_descriptor m_t4;
    // Enables sequence termination when coverage goals are met
    bit m_terminateOnCoverageGoalsMet = 1;
    // Enables sequence termination when distribution replay data ends
    bit m_terminateOnReplayEnd = 1;
    bit m_replayEndReached = 0;
    // Enables sequence termination after a specific number of sequence items
    int m_iterationLimit = 0;
    // Tracks number of iterations
    int m_iterationCount = 0;
    // Controls how often a coverage report is produced
    int m_coverageReportInterval = 1;
    longint                              m_t1__ll_desc_tot_sz__size;
    longint                              m_t1__ll_desc_tot_sz__sum;
    longint                              m_t2__ll_desc_tot_sz__size;
    longint                              m_t2__ll_desc_tot_sz__sum;
    longint                              m_t3__ll_desc_tot_sz__size;
    longint                              m_t3__ll_desc_tot_sz__sum;
    longint                              m_t4__ll_desc_tot_sz__size;
    longint                              m_t4__ll_desc_tot_sz__sum;


// Coverage Strategy fields
    wb_dma_infact_4par_sw_seq_pc_closure #(wb_dma_infact_4par_sw_seq_t)       m_pc_closure;

//</item_fields>
    
//<user_data,gen>

//</user_data>
     

    //***************************************************************
    //* new()
    //***************************************************************
    function new(string name="");
    	super.new(name);
    endfunction
    
    //***************************************************************
    //* body()
    //***************************************************************
    virtual task body();
    	// Create the inFact scheduler
    	m_scheduler = new(get_full_name());
    	
    	// Register action tasks with the scheduler
    	register_actions();
    
        // Create Coverage Strategies
        create_cov_strategies();
    
    	// Run all the test engines
    	m_scheduler.run_all();
    	
    	// Clean up after the test engines return
//<delete_testengines,gen>
        begin
            inFactSv::TestEngine   te;
            te = m_scheduler.wb_dma_infact_4par_sw_seq();
            te.delete();

        end
//</delete_testengines>
    	
    endtask
    
    
    //***************************************************************
    //* Action Tasks
    //***************************************************************
//<action_tasks>

//<action::_infact_checkcov::()>
    //***************************************************************
    //* Action task action_infact_checkcov
    //* Displays coverage report 

    //**************************************************************** 
   virtual task action_infact_checkcov();
        begin
            bit ending = 0;
            m_iterationCount++;
            if ((m_iterationLimit > 0 && 
                m_iterationCount >= m_iterationLimit) ||
                (m_terminateOnCoverageGoalsMet && allCoverageGoalsHaveBeenMet())) begin
                ending = 1;
            end
            // Display a coverage report when requested or when the sequence ends
            if (m_coverageReportInterval > 0 && 
                (ending || !(m_iterationCount % m_coverageReportInterval))) begin
                string report = getCoverageReport();
                if (report != "") begin
                    `uvm_info(get_full_name(), {"Coverage Report:\n", report}, UVM_MEDIUM);
                end
            end
            if (m_terminateOnReplayEnd && m_replayEndReached) begin
      `uvm_info(get_full_name(), "Reached end of replay data. Ending sequence", UVM_MEDIUM);
      ending = 1;
    end
    if (ending) begin
                m_te.stop_loop_expansion_after(0, m_te.loop_depth()-1);
            end
        end

    endtask
//</action::_infact_checkcov::()>


























































































































































































































































































































































































































































//<action::_init_xfer__t4__end::()>
    //***************************************************************
    //* Action task action_init_xfer__t4__end
    //**************************************************************** 
   virtual task action_init_xfer__t4__end();
                if (m_terminateOnReplayEnd && m_replayEndReached) begin
          `uvm_info(get_full_name(), "Skipping finish_item due to replay end", UVM_MEDIUM);
        end else begin
          finish_item(m_t4);
        end

    endtask
//</action::_init_xfer__t4__end::()>

//<action::_init_xfer__t4__begin::()>
    //***************************************************************
    //* Action task action_init_xfer__t4__begin
    //**************************************************************** 
   virtual task action_init_xfer__t4__begin();
        m_t4 = wb_dma_descriptor::type_id::create();
        if (m_terminateOnReplayEnd && m_replayEndReached) begin
          `uvm_info(get_full_name(), "Skipping start_item due to replay end", UVM_MEDIUM);
        end else begin
          start_item(m_t4);
        end

    endtask
//</action::_init_xfer__t4__begin::()>

//<action::_init_xfer__t3__end::()>
    //***************************************************************
    //* Action task action_init_xfer__t3__end
    //**************************************************************** 
   virtual task action_init_xfer__t3__end();
                if (m_terminateOnReplayEnd && m_replayEndReached) begin
          `uvm_info(get_full_name(), "Skipping finish_item due to replay end", UVM_MEDIUM);
        end else begin
          finish_item(m_t3);
        end

    endtask
//</action::_init_xfer__t3__end::()>

//<action::_init_xfer__t3__begin::()>
    //***************************************************************
    //* Action task action_init_xfer__t3__begin
    //**************************************************************** 
   virtual task action_init_xfer__t3__begin();
        m_t3 = wb_dma_descriptor::type_id::create();
        if (m_terminateOnReplayEnd && m_replayEndReached) begin
          `uvm_info(get_full_name(), "Skipping start_item due to replay end", UVM_MEDIUM);
        end else begin
          start_item(m_t3);
        end

    endtask
//</action::_init_xfer__t3__begin::()>

//<action::_init_xfer__t2__end::()>
    //***************************************************************
    //* Action task action_init_xfer__t2__end
    //**************************************************************** 
   virtual task action_init_xfer__t2__end();
                if (m_terminateOnReplayEnd && m_replayEndReached) begin
          `uvm_info(get_full_name(), "Skipping finish_item due to replay end", UVM_MEDIUM);
        end else begin
          finish_item(m_t2);
        end

    endtask
//</action::_init_xfer__t2__end::()>

//<action::_init_xfer__t2__begin::()>
    //***************************************************************
    //* Action task action_init_xfer__t2__begin
    //**************************************************************** 
   virtual task action_init_xfer__t2__begin();
        m_t2 = wb_dma_descriptor::type_id::create();
        if (m_terminateOnReplayEnd && m_replayEndReached) begin
          `uvm_info(get_full_name(), "Skipping start_item due to replay end", UVM_MEDIUM);
        end else begin
          start_item(m_t2);
        end

    endtask
//</action::_init_xfer__t2__begin::()>

//<action::_init_xfer__t1__end::()>
    //***************************************************************
    //* Action task action_init_xfer__t1__end
    //**************************************************************** 
   virtual task action_init_xfer__t1__end();
                if (m_terminateOnReplayEnd && m_replayEndReached) begin
          `uvm_info(get_full_name(), "Skipping finish_item due to replay end", UVM_MEDIUM);
        end else begin
          finish_item(m_t1);
        end

    endtask
//</action::_init_xfer__t1__end::()>

//<action::_init_xfer__t1__begin::()>
    //***************************************************************
    //* Action task action_init_xfer__t1__begin
    //**************************************************************** 
   virtual task action_init_xfer__t1__begin();
        m_t1 = wb_dma_descriptor::type_id::create();
        if (m_terminateOnReplayEnd && m_replayEndReached) begin
          `uvm_info(get_full_name(), "Skipping start_item due to replay end", UVM_MEDIUM);
        end else begin
          start_item(m_t1);
        end

    endtask
//</action::_init_xfer__t1__begin::()>

//<action::_init::(##a15a1c9061d180c45065bc9fc24cf98e)>
    //***************************************************************
    //* Action task action_init
    //* action_stmt = m_iterationLimit = 16;
    //**************************************************************** 
   virtual task action_init();
        m_iterationLimit = 16;
    endtask
//</action::_init::(##a15a1c9061d180c45065bc9fc24cf98e)>

//<signed_meta_action::_t4__ll_desc_tot_sz__sum::()>
    //***************************************************************
    //* Action task action_t4__ll_desc_tot_sz__sum
    //**************************************************************** 
   virtual task action_t4__ll_desc_tot_sz__sum(longint meta_val);
        m_t4__ll_desc_tot_sz__sum = meta_val;
    endtask
//</signed_meta_action::_t4__ll_desc_tot_sz__sum::()>

//<signed_meta_action::_t3__ll_desc_tot_sz__sum::()>
    //***************************************************************
    //* Action task action_t3__ll_desc_tot_sz__sum
    //**************************************************************** 
   virtual task action_t3__ll_desc_tot_sz__sum(longint meta_val);
        m_t3__ll_desc_tot_sz__sum = meta_val;
    endtask
//</signed_meta_action::_t3__ll_desc_tot_sz__sum::()>

//<signed_meta_action::_t2__ll_desc_tot_sz__sum::()>
    //***************************************************************
    //* Action task action_t2__ll_desc_tot_sz__sum
    //**************************************************************** 
   virtual task action_t2__ll_desc_tot_sz__sum(longint meta_val);
        m_t2__ll_desc_tot_sz__sum = meta_val;
    endtask
//</signed_meta_action::_t2__ll_desc_tot_sz__sum::()>

//<signed_meta_action::_t1__ll_desc_tot_sz__sum::()>
    //***************************************************************
    //* Action task action_t1__ll_desc_tot_sz__sum
    //**************************************************************** 
   virtual task action_t1__ll_desc_tot_sz__sum(longint meta_val);
        m_t1__ll_desc_tot_sz__sum = meta_val;
    endtask
//</signed_meta_action::_t1__ll_desc_tot_sz__sum::()>

//<unsigned_meta_action::_t4__transfer_sz::()>
    //***************************************************************
    //* Action task action_t4__transfer_sz
    //**************************************************************** 
   virtual task action_t4__transfer_sz(longint unsigned meta_val);
        m_t4.transfer_sz = meta_val;
    endtask
//</unsigned_meta_action::_t4__transfer_sz::()>

//<unsigned_meta_action::_t4__ll_desc_tot_sz__15__::()>
    //***************************************************************
    //* Action task action_t4__ll_desc_tot_sz__15__
    //**************************************************************** 
   virtual task action_t4__ll_desc_tot_sz__15__(longint unsigned meta_val);
        m_t4.ll_desc_tot_sz[15] = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc_tot_sz__15__::()>

//<unsigned_meta_action::_t4__ll_desc_tot_sz__14__::()>
    //***************************************************************
    //* Action task action_t4__ll_desc_tot_sz__14__
    //**************************************************************** 
   virtual task action_t4__ll_desc_tot_sz__14__(longint unsigned meta_val);
        m_t4.ll_desc_tot_sz[14] = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc_tot_sz__14__::()>

//<unsigned_meta_action::_t4__ll_desc_tot_sz__13__::()>
    //***************************************************************
    //* Action task action_t4__ll_desc_tot_sz__13__
    //**************************************************************** 
   virtual task action_t4__ll_desc_tot_sz__13__(longint unsigned meta_val);
        m_t4.ll_desc_tot_sz[13] = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc_tot_sz__13__::()>

//<unsigned_meta_action::_t4__ll_desc_tot_sz__12__::()>
    //***************************************************************
    //* Action task action_t4__ll_desc_tot_sz__12__
    //**************************************************************** 
   virtual task action_t4__ll_desc_tot_sz__12__(longint unsigned meta_val);
        m_t4.ll_desc_tot_sz[12] = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc_tot_sz__12__::()>

//<unsigned_meta_action::_t4__ll_desc_tot_sz__11__::()>
    //***************************************************************
    //* Action task action_t4__ll_desc_tot_sz__11__
    //**************************************************************** 
   virtual task action_t4__ll_desc_tot_sz__11__(longint unsigned meta_val);
        m_t4.ll_desc_tot_sz[11] = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc_tot_sz__11__::()>

//<unsigned_meta_action::_t4__ll_desc_tot_sz__10__::()>
    //***************************************************************
    //* Action task action_t4__ll_desc_tot_sz__10__
    //**************************************************************** 
   virtual task action_t4__ll_desc_tot_sz__10__(longint unsigned meta_val);
        m_t4.ll_desc_tot_sz[10] = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc_tot_sz__10__::()>

//<unsigned_meta_action::_t4__ll_desc_tot_sz__9__::()>
    //***************************************************************
    //* Action task action_t4__ll_desc_tot_sz__9__
    //**************************************************************** 
   virtual task action_t4__ll_desc_tot_sz__9__(longint unsigned meta_val);
        m_t4.ll_desc_tot_sz[9] = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc_tot_sz__9__::()>

//<unsigned_meta_action::_t4__ll_desc_tot_sz__8__::()>
    //***************************************************************
    //* Action task action_t4__ll_desc_tot_sz__8__
    //**************************************************************** 
   virtual task action_t4__ll_desc_tot_sz__8__(longint unsigned meta_val);
        m_t4.ll_desc_tot_sz[8] = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc_tot_sz__8__::()>

//<unsigned_meta_action::_t4__ll_desc_tot_sz__7__::()>
    //***************************************************************
    //* Action task action_t4__ll_desc_tot_sz__7__
    //**************************************************************** 
   virtual task action_t4__ll_desc_tot_sz__7__(longint unsigned meta_val);
        m_t4.ll_desc_tot_sz[7] = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc_tot_sz__7__::()>

//<unsigned_meta_action::_t4__ll_desc_tot_sz__6__::()>
    //***************************************************************
    //* Action task action_t4__ll_desc_tot_sz__6__
    //**************************************************************** 
   virtual task action_t4__ll_desc_tot_sz__6__(longint unsigned meta_val);
        m_t4.ll_desc_tot_sz[6] = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc_tot_sz__6__::()>

//<unsigned_meta_action::_t4__ll_desc_tot_sz__5__::()>
    //***************************************************************
    //* Action task action_t4__ll_desc_tot_sz__5__
    //**************************************************************** 
   virtual task action_t4__ll_desc_tot_sz__5__(longint unsigned meta_val);
        m_t4.ll_desc_tot_sz[5] = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc_tot_sz__5__::()>

//<unsigned_meta_action::_t4__ll_desc_tot_sz__4__::()>
    //***************************************************************
    //* Action task action_t4__ll_desc_tot_sz__4__
    //**************************************************************** 
   virtual task action_t4__ll_desc_tot_sz__4__(longint unsigned meta_val);
        m_t4.ll_desc_tot_sz[4] = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc_tot_sz__4__::()>

//<unsigned_meta_action::_t4__ll_desc_tot_sz__3__::()>
    //***************************************************************
    //* Action task action_t4__ll_desc_tot_sz__3__
    //**************************************************************** 
   virtual task action_t4__ll_desc_tot_sz__3__(longint unsigned meta_val);
        m_t4.ll_desc_tot_sz[3] = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc_tot_sz__3__::()>

//<unsigned_meta_action::_t4__ll_desc_tot_sz__2__::()>
    //***************************************************************
    //* Action task action_t4__ll_desc_tot_sz__2__
    //**************************************************************** 
   virtual task action_t4__ll_desc_tot_sz__2__(longint unsigned meta_val);
        m_t4.ll_desc_tot_sz[2] = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc_tot_sz__2__::()>

//<unsigned_meta_action::_t4__ll_desc_tot_sz__1__::()>
    //***************************************************************
    //* Action task action_t4__ll_desc_tot_sz__1__
    //**************************************************************** 
   virtual task action_t4__ll_desc_tot_sz__1__(longint unsigned meta_val);
        m_t4.ll_desc_tot_sz[1] = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc_tot_sz__1__::()>

//<unsigned_meta_action::_t4__ll_desc_tot_sz__0__::()>
    //***************************************************************
    //* Action task action_t4__ll_desc_tot_sz__0__
    //**************************************************************** 
   virtual task action_t4__ll_desc_tot_sz__0__(longint unsigned meta_val);
        m_t4.ll_desc_tot_sz[0] = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc_tot_sz__0__::()>

//<unsigned_meta_action::_t4__ll_desc_sz::()>
    //***************************************************************
    //* Action task action_t4__ll_desc_sz
    //**************************************************************** 
   virtual task action_t4__ll_desc_sz(longint unsigned meta_val);
        m_t4.ll_desc_sz = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc_sz::()>

//<unsigned_meta_action::_t4__ll_desc__15____tot_sz::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__15____tot_sz
    //**************************************************************** 
   virtual task action_t4__ll_desc__15____tot_sz(longint unsigned meta_val);
        m_t4.ll_desc[15].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__15____tot_sz::()>

//<unsigned_meta_action::_t4__ll_desc__15____dst_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__15____dst_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__15____dst_sel(longint unsigned meta_val);
        m_t4.ll_desc[15].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__15____dst_sel::()>

//<unsigned_meta_action::_t4__ll_desc__15____src_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__15____src_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__15____src_sel(longint unsigned meta_val);
        m_t4.ll_desc[15].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__15____src_sel::()>

//<unsigned_meta_action::_t4__ll_desc__15____inc_dst::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__15____inc_dst
    //**************************************************************** 
   virtual task action_t4__ll_desc__15____inc_dst(longint unsigned meta_val);
        m_t4.ll_desc[15].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__15____inc_dst::()>

//<unsigned_meta_action::_t4__ll_desc__15____inc_src::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__15____inc_src
    //**************************************************************** 
   virtual task action_t4__ll_desc__15____inc_src(longint unsigned meta_val);
        m_t4.ll_desc[15].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__15____inc_src::()>

//<unsigned_meta_action::_t4__ll_desc__14____tot_sz::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__14____tot_sz
    //**************************************************************** 
   virtual task action_t4__ll_desc__14____tot_sz(longint unsigned meta_val);
        m_t4.ll_desc[14].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__14____tot_sz::()>

//<unsigned_meta_action::_t4__ll_desc__14____dst_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__14____dst_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__14____dst_sel(longint unsigned meta_val);
        m_t4.ll_desc[14].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__14____dst_sel::()>

//<unsigned_meta_action::_t4__ll_desc__14____src_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__14____src_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__14____src_sel(longint unsigned meta_val);
        m_t4.ll_desc[14].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__14____src_sel::()>

//<unsigned_meta_action::_t4__ll_desc__14____inc_dst::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__14____inc_dst
    //**************************************************************** 
   virtual task action_t4__ll_desc__14____inc_dst(longint unsigned meta_val);
        m_t4.ll_desc[14].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__14____inc_dst::()>

//<unsigned_meta_action::_t4__ll_desc__14____inc_src::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__14____inc_src
    //**************************************************************** 
   virtual task action_t4__ll_desc__14____inc_src(longint unsigned meta_val);
        m_t4.ll_desc[14].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__14____inc_src::()>

//<unsigned_meta_action::_t4__ll_desc__13____tot_sz::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__13____tot_sz
    //**************************************************************** 
   virtual task action_t4__ll_desc__13____tot_sz(longint unsigned meta_val);
        m_t4.ll_desc[13].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__13____tot_sz::()>

//<unsigned_meta_action::_t4__ll_desc__13____dst_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__13____dst_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__13____dst_sel(longint unsigned meta_val);
        m_t4.ll_desc[13].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__13____dst_sel::()>

//<unsigned_meta_action::_t4__ll_desc__13____src_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__13____src_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__13____src_sel(longint unsigned meta_val);
        m_t4.ll_desc[13].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__13____src_sel::()>

//<unsigned_meta_action::_t4__ll_desc__13____inc_dst::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__13____inc_dst
    //**************************************************************** 
   virtual task action_t4__ll_desc__13____inc_dst(longint unsigned meta_val);
        m_t4.ll_desc[13].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__13____inc_dst::()>

//<unsigned_meta_action::_t4__ll_desc__13____inc_src::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__13____inc_src
    //**************************************************************** 
   virtual task action_t4__ll_desc__13____inc_src(longint unsigned meta_val);
        m_t4.ll_desc[13].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__13____inc_src::()>

//<unsigned_meta_action::_t4__ll_desc__12____tot_sz::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__12____tot_sz
    //**************************************************************** 
   virtual task action_t4__ll_desc__12____tot_sz(longint unsigned meta_val);
        m_t4.ll_desc[12].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__12____tot_sz::()>

//<unsigned_meta_action::_t4__ll_desc__12____dst_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__12____dst_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__12____dst_sel(longint unsigned meta_val);
        m_t4.ll_desc[12].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__12____dst_sel::()>

//<unsigned_meta_action::_t4__ll_desc__12____src_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__12____src_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__12____src_sel(longint unsigned meta_val);
        m_t4.ll_desc[12].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__12____src_sel::()>

//<unsigned_meta_action::_t4__ll_desc__12____inc_dst::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__12____inc_dst
    //**************************************************************** 
   virtual task action_t4__ll_desc__12____inc_dst(longint unsigned meta_val);
        m_t4.ll_desc[12].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__12____inc_dst::()>

//<unsigned_meta_action::_t4__ll_desc__12____inc_src::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__12____inc_src
    //**************************************************************** 
   virtual task action_t4__ll_desc__12____inc_src(longint unsigned meta_val);
        m_t4.ll_desc[12].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__12____inc_src::()>

//<unsigned_meta_action::_t4__ll_desc__11____tot_sz::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__11____tot_sz
    //**************************************************************** 
   virtual task action_t4__ll_desc__11____tot_sz(longint unsigned meta_val);
        m_t4.ll_desc[11].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__11____tot_sz::()>

//<unsigned_meta_action::_t4__ll_desc__11____dst_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__11____dst_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__11____dst_sel(longint unsigned meta_val);
        m_t4.ll_desc[11].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__11____dst_sel::()>

//<unsigned_meta_action::_t4__ll_desc__11____src_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__11____src_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__11____src_sel(longint unsigned meta_val);
        m_t4.ll_desc[11].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__11____src_sel::()>

//<unsigned_meta_action::_t4__ll_desc__11____inc_dst::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__11____inc_dst
    //**************************************************************** 
   virtual task action_t4__ll_desc__11____inc_dst(longint unsigned meta_val);
        m_t4.ll_desc[11].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__11____inc_dst::()>

//<unsigned_meta_action::_t4__ll_desc__11____inc_src::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__11____inc_src
    //**************************************************************** 
   virtual task action_t4__ll_desc__11____inc_src(longint unsigned meta_val);
        m_t4.ll_desc[11].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__11____inc_src::()>

//<unsigned_meta_action::_t4__ll_desc__10____tot_sz::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__10____tot_sz
    //**************************************************************** 
   virtual task action_t4__ll_desc__10____tot_sz(longint unsigned meta_val);
        m_t4.ll_desc[10].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__10____tot_sz::()>

//<unsigned_meta_action::_t4__ll_desc__10____dst_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__10____dst_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__10____dst_sel(longint unsigned meta_val);
        m_t4.ll_desc[10].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__10____dst_sel::()>

//<unsigned_meta_action::_t4__ll_desc__10____src_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__10____src_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__10____src_sel(longint unsigned meta_val);
        m_t4.ll_desc[10].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__10____src_sel::()>

//<unsigned_meta_action::_t4__ll_desc__10____inc_dst::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__10____inc_dst
    //**************************************************************** 
   virtual task action_t4__ll_desc__10____inc_dst(longint unsigned meta_val);
        m_t4.ll_desc[10].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__10____inc_dst::()>

//<unsigned_meta_action::_t4__ll_desc__10____inc_src::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__10____inc_src
    //**************************************************************** 
   virtual task action_t4__ll_desc__10____inc_src(longint unsigned meta_val);
        m_t4.ll_desc[10].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__10____inc_src::()>

//<unsigned_meta_action::_t4__ll_desc__9____tot_sz::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__9____tot_sz
    //**************************************************************** 
   virtual task action_t4__ll_desc__9____tot_sz(longint unsigned meta_val);
        m_t4.ll_desc[9].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__9____tot_sz::()>

//<unsigned_meta_action::_t4__ll_desc__9____dst_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__9____dst_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__9____dst_sel(longint unsigned meta_val);
        m_t4.ll_desc[9].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__9____dst_sel::()>

//<unsigned_meta_action::_t4__ll_desc__9____src_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__9____src_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__9____src_sel(longint unsigned meta_val);
        m_t4.ll_desc[9].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__9____src_sel::()>

//<unsigned_meta_action::_t4__ll_desc__9____inc_dst::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__9____inc_dst
    //**************************************************************** 
   virtual task action_t4__ll_desc__9____inc_dst(longint unsigned meta_val);
        m_t4.ll_desc[9].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__9____inc_dst::()>

//<unsigned_meta_action::_t4__ll_desc__9____inc_src::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__9____inc_src
    //**************************************************************** 
   virtual task action_t4__ll_desc__9____inc_src(longint unsigned meta_val);
        m_t4.ll_desc[9].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__9____inc_src::()>

//<unsigned_meta_action::_t4__ll_desc__8____tot_sz::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__8____tot_sz
    //**************************************************************** 
   virtual task action_t4__ll_desc__8____tot_sz(longint unsigned meta_val);
        m_t4.ll_desc[8].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__8____tot_sz::()>

//<unsigned_meta_action::_t4__ll_desc__8____dst_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__8____dst_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__8____dst_sel(longint unsigned meta_val);
        m_t4.ll_desc[8].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__8____dst_sel::()>

//<unsigned_meta_action::_t4__ll_desc__8____src_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__8____src_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__8____src_sel(longint unsigned meta_val);
        m_t4.ll_desc[8].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__8____src_sel::()>

//<unsigned_meta_action::_t4__ll_desc__8____inc_dst::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__8____inc_dst
    //**************************************************************** 
   virtual task action_t4__ll_desc__8____inc_dst(longint unsigned meta_val);
        m_t4.ll_desc[8].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__8____inc_dst::()>

//<unsigned_meta_action::_t4__ll_desc__8____inc_src::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__8____inc_src
    //**************************************************************** 
   virtual task action_t4__ll_desc__8____inc_src(longint unsigned meta_val);
        m_t4.ll_desc[8].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__8____inc_src::()>

//<unsigned_meta_action::_t4__ll_desc__7____tot_sz::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__7____tot_sz
    //**************************************************************** 
   virtual task action_t4__ll_desc__7____tot_sz(longint unsigned meta_val);
        m_t4.ll_desc[7].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__7____tot_sz::()>

//<unsigned_meta_action::_t4__ll_desc__7____dst_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__7____dst_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__7____dst_sel(longint unsigned meta_val);
        m_t4.ll_desc[7].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__7____dst_sel::()>

//<unsigned_meta_action::_t4__ll_desc__7____src_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__7____src_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__7____src_sel(longint unsigned meta_val);
        m_t4.ll_desc[7].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__7____src_sel::()>

//<unsigned_meta_action::_t4__ll_desc__7____inc_dst::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__7____inc_dst
    //**************************************************************** 
   virtual task action_t4__ll_desc__7____inc_dst(longint unsigned meta_val);
        m_t4.ll_desc[7].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__7____inc_dst::()>

//<unsigned_meta_action::_t4__ll_desc__7____inc_src::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__7____inc_src
    //**************************************************************** 
   virtual task action_t4__ll_desc__7____inc_src(longint unsigned meta_val);
        m_t4.ll_desc[7].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__7____inc_src::()>

//<unsigned_meta_action::_t4__ll_desc__6____tot_sz::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__6____tot_sz
    //**************************************************************** 
   virtual task action_t4__ll_desc__6____tot_sz(longint unsigned meta_val);
        m_t4.ll_desc[6].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__6____tot_sz::()>

//<unsigned_meta_action::_t4__ll_desc__6____dst_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__6____dst_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__6____dst_sel(longint unsigned meta_val);
        m_t4.ll_desc[6].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__6____dst_sel::()>

//<unsigned_meta_action::_t4__ll_desc__6____src_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__6____src_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__6____src_sel(longint unsigned meta_val);
        m_t4.ll_desc[6].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__6____src_sel::()>

//<unsigned_meta_action::_t4__ll_desc__6____inc_dst::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__6____inc_dst
    //**************************************************************** 
   virtual task action_t4__ll_desc__6____inc_dst(longint unsigned meta_val);
        m_t4.ll_desc[6].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__6____inc_dst::()>

//<unsigned_meta_action::_t4__ll_desc__6____inc_src::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__6____inc_src
    //**************************************************************** 
   virtual task action_t4__ll_desc__6____inc_src(longint unsigned meta_val);
        m_t4.ll_desc[6].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__6____inc_src::()>

//<unsigned_meta_action::_t4__ll_desc__5____tot_sz::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__5____tot_sz
    //**************************************************************** 
   virtual task action_t4__ll_desc__5____tot_sz(longint unsigned meta_val);
        m_t4.ll_desc[5].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__5____tot_sz::()>

//<unsigned_meta_action::_t4__ll_desc__5____dst_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__5____dst_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__5____dst_sel(longint unsigned meta_val);
        m_t4.ll_desc[5].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__5____dst_sel::()>

//<unsigned_meta_action::_t4__ll_desc__5____src_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__5____src_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__5____src_sel(longint unsigned meta_val);
        m_t4.ll_desc[5].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__5____src_sel::()>

//<unsigned_meta_action::_t4__ll_desc__5____inc_dst::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__5____inc_dst
    //**************************************************************** 
   virtual task action_t4__ll_desc__5____inc_dst(longint unsigned meta_val);
        m_t4.ll_desc[5].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__5____inc_dst::()>

//<unsigned_meta_action::_t4__ll_desc__5____inc_src::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__5____inc_src
    //**************************************************************** 
   virtual task action_t4__ll_desc__5____inc_src(longint unsigned meta_val);
        m_t4.ll_desc[5].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__5____inc_src::()>

//<unsigned_meta_action::_t4__ll_desc__4____tot_sz::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__4____tot_sz
    //**************************************************************** 
   virtual task action_t4__ll_desc__4____tot_sz(longint unsigned meta_val);
        m_t4.ll_desc[4].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__4____tot_sz::()>

//<unsigned_meta_action::_t4__ll_desc__4____dst_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__4____dst_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__4____dst_sel(longint unsigned meta_val);
        m_t4.ll_desc[4].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__4____dst_sel::()>

//<unsigned_meta_action::_t4__ll_desc__4____src_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__4____src_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__4____src_sel(longint unsigned meta_val);
        m_t4.ll_desc[4].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__4____src_sel::()>

//<unsigned_meta_action::_t4__ll_desc__4____inc_dst::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__4____inc_dst
    //**************************************************************** 
   virtual task action_t4__ll_desc__4____inc_dst(longint unsigned meta_val);
        m_t4.ll_desc[4].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__4____inc_dst::()>

//<unsigned_meta_action::_t4__ll_desc__4____inc_src::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__4____inc_src
    //**************************************************************** 
   virtual task action_t4__ll_desc__4____inc_src(longint unsigned meta_val);
        m_t4.ll_desc[4].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__4____inc_src::()>

//<unsigned_meta_action::_t4__ll_desc__3____tot_sz::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__3____tot_sz
    //**************************************************************** 
   virtual task action_t4__ll_desc__3____tot_sz(longint unsigned meta_val);
        m_t4.ll_desc[3].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__3____tot_sz::()>

//<unsigned_meta_action::_t4__ll_desc__3____dst_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__3____dst_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__3____dst_sel(longint unsigned meta_val);
        m_t4.ll_desc[3].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__3____dst_sel::()>

//<unsigned_meta_action::_t4__ll_desc__3____src_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__3____src_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__3____src_sel(longint unsigned meta_val);
        m_t4.ll_desc[3].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__3____src_sel::()>

//<unsigned_meta_action::_t4__ll_desc__3____inc_dst::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__3____inc_dst
    //**************************************************************** 
   virtual task action_t4__ll_desc__3____inc_dst(longint unsigned meta_val);
        m_t4.ll_desc[3].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__3____inc_dst::()>

//<unsigned_meta_action::_t4__ll_desc__3____inc_src::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__3____inc_src
    //**************************************************************** 
   virtual task action_t4__ll_desc__3____inc_src(longint unsigned meta_val);
        m_t4.ll_desc[3].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__3____inc_src::()>

//<unsigned_meta_action::_t4__ll_desc__2____tot_sz::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__2____tot_sz
    //**************************************************************** 
   virtual task action_t4__ll_desc__2____tot_sz(longint unsigned meta_val);
        m_t4.ll_desc[2].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__2____tot_sz::()>

//<unsigned_meta_action::_t4__ll_desc__2____dst_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__2____dst_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__2____dst_sel(longint unsigned meta_val);
        m_t4.ll_desc[2].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__2____dst_sel::()>

//<unsigned_meta_action::_t4__ll_desc__2____src_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__2____src_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__2____src_sel(longint unsigned meta_val);
        m_t4.ll_desc[2].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__2____src_sel::()>

//<unsigned_meta_action::_t4__ll_desc__2____inc_dst::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__2____inc_dst
    //**************************************************************** 
   virtual task action_t4__ll_desc__2____inc_dst(longint unsigned meta_val);
        m_t4.ll_desc[2].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__2____inc_dst::()>

//<unsigned_meta_action::_t4__ll_desc__2____inc_src::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__2____inc_src
    //**************************************************************** 
   virtual task action_t4__ll_desc__2____inc_src(longint unsigned meta_val);
        m_t4.ll_desc[2].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__2____inc_src::()>

//<unsigned_meta_action::_t4__ll_desc__1____tot_sz::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__1____tot_sz
    //**************************************************************** 
   virtual task action_t4__ll_desc__1____tot_sz(longint unsigned meta_val);
        m_t4.ll_desc[1].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__1____tot_sz::()>

//<unsigned_meta_action::_t4__ll_desc__1____dst_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__1____dst_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__1____dst_sel(longint unsigned meta_val);
        m_t4.ll_desc[1].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__1____dst_sel::()>

//<unsigned_meta_action::_t4__ll_desc__1____src_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__1____src_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__1____src_sel(longint unsigned meta_val);
        m_t4.ll_desc[1].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__1____src_sel::()>

//<unsigned_meta_action::_t4__ll_desc__1____inc_dst::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__1____inc_dst
    //**************************************************************** 
   virtual task action_t4__ll_desc__1____inc_dst(longint unsigned meta_val);
        m_t4.ll_desc[1].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__1____inc_dst::()>

//<unsigned_meta_action::_t4__ll_desc__1____inc_src::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__1____inc_src
    //**************************************************************** 
   virtual task action_t4__ll_desc__1____inc_src(longint unsigned meta_val);
        m_t4.ll_desc[1].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__1____inc_src::()>

//<unsigned_meta_action::_t4__ll_desc__0____tot_sz::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__0____tot_sz
    //**************************************************************** 
   virtual task action_t4__ll_desc__0____tot_sz(longint unsigned meta_val);
        m_t4.ll_desc[0].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__0____tot_sz::()>

//<unsigned_meta_action::_t4__ll_desc__0____dst_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__0____dst_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__0____dst_sel(longint unsigned meta_val);
        m_t4.ll_desc[0].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__0____dst_sel::()>

//<unsigned_meta_action::_t4__ll_desc__0____src_sel::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__0____src_sel
    //**************************************************************** 
   virtual task action_t4__ll_desc__0____src_sel(longint unsigned meta_val);
        m_t4.ll_desc[0].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__0____src_sel::()>

//<unsigned_meta_action::_t4__ll_desc__0____inc_dst::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__0____inc_dst
    //**************************************************************** 
   virtual task action_t4__ll_desc__0____inc_dst(longint unsigned meta_val);
        m_t4.ll_desc[0].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__0____inc_dst::()>

//<unsigned_meta_action::_t4__ll_desc__0____inc_src::()>
    //***************************************************************
    //* Action task action_t4__ll_desc__0____inc_src
    //**************************************************************** 
   virtual task action_t4__ll_desc__0____inc_src(longint unsigned meta_val);
        m_t4.ll_desc[0].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t4__ll_desc__0____inc_src::()>

//<unsigned_meta_action::_t4__chk_sz::()>
    //***************************************************************
    //* Action task action_t4__chk_sz
    //**************************************************************** 
   virtual task action_t4__chk_sz(longint unsigned meta_val);
        m_t4.chk_sz = meta_val;
    endtask
//</unsigned_meta_action::_t4__chk_sz::()>

//<unsigned_meta_action::_t4__tot_sz::()>
    //***************************************************************
    //* Action task action_t4__tot_sz
    //**************************************************************** 
   virtual task action_t4__tot_sz(longint unsigned meta_val);
        m_t4.tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t4__tot_sz::()>

//<unsigned_meta_action::_t4__dst_sel::()>
    //***************************************************************
    //* Action task action_t4__dst_sel
    //**************************************************************** 
   virtual task action_t4__dst_sel(longint unsigned meta_val);
        m_t4.dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__dst_sel::()>

//<unsigned_meta_action::_t4__src_sel::()>
    //***************************************************************
    //* Action task action_t4__src_sel
    //**************************************************************** 
   virtual task action_t4__src_sel(longint unsigned meta_val);
        m_t4.src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t4__src_sel::()>

//<unsigned_meta_action::_t4__inc_dst::()>
    //***************************************************************
    //* Action task action_t4__inc_dst
    //**************************************************************** 
   virtual task action_t4__inc_dst(longint unsigned meta_val);
        m_t4.inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t4__inc_dst::()>

//<unsigned_meta_action::_t4__inc_src::()>
    //***************************************************************
    //* Action task action_t4__inc_src
    //**************************************************************** 
   virtual task action_t4__inc_src(longint unsigned meta_val);
        m_t4.inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t4__inc_src::()>

//<unsigned_meta_action::_t4__mode::()>
    //***************************************************************
    //* Action task action_t4__mode
    //**************************************************************** 
   virtual task action_t4__mode(longint unsigned meta_val);
        m_t4.mode = meta_val;
    endtask
//</unsigned_meta_action::_t4__mode::()>

//<unsigned_meta_action::_t4__channel::()>
    //***************************************************************
    //* Action task action_t4__channel
    //**************************************************************** 
   virtual task action_t4__channel(longint unsigned meta_val);
        m_t4.channel = meta_val;
    endtask
//</unsigned_meta_action::_t4__channel::()>

//<unsigned_meta_action::_t3__transfer_sz::()>
    //***************************************************************
    //* Action task action_t3__transfer_sz
    //**************************************************************** 
   virtual task action_t3__transfer_sz(longint unsigned meta_val);
        m_t3.transfer_sz = meta_val;
    endtask
//</unsigned_meta_action::_t3__transfer_sz::()>

//<unsigned_meta_action::_t3__ll_desc_tot_sz__15__::()>
    //***************************************************************
    //* Action task action_t3__ll_desc_tot_sz__15__
    //**************************************************************** 
   virtual task action_t3__ll_desc_tot_sz__15__(longint unsigned meta_val);
        m_t3.ll_desc_tot_sz[15] = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc_tot_sz__15__::()>

//<unsigned_meta_action::_t3__ll_desc_tot_sz__14__::()>
    //***************************************************************
    //* Action task action_t3__ll_desc_tot_sz__14__
    //**************************************************************** 
   virtual task action_t3__ll_desc_tot_sz__14__(longint unsigned meta_val);
        m_t3.ll_desc_tot_sz[14] = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc_tot_sz__14__::()>

//<unsigned_meta_action::_t3__ll_desc_tot_sz__13__::()>
    //***************************************************************
    //* Action task action_t3__ll_desc_tot_sz__13__
    //**************************************************************** 
   virtual task action_t3__ll_desc_tot_sz__13__(longint unsigned meta_val);
        m_t3.ll_desc_tot_sz[13] = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc_tot_sz__13__::()>

//<unsigned_meta_action::_t3__ll_desc_tot_sz__12__::()>
    //***************************************************************
    //* Action task action_t3__ll_desc_tot_sz__12__
    //**************************************************************** 
   virtual task action_t3__ll_desc_tot_sz__12__(longint unsigned meta_val);
        m_t3.ll_desc_tot_sz[12] = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc_tot_sz__12__::()>

//<unsigned_meta_action::_t3__ll_desc_tot_sz__11__::()>
    //***************************************************************
    //* Action task action_t3__ll_desc_tot_sz__11__
    //**************************************************************** 
   virtual task action_t3__ll_desc_tot_sz__11__(longint unsigned meta_val);
        m_t3.ll_desc_tot_sz[11] = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc_tot_sz__11__::()>

//<unsigned_meta_action::_t3__ll_desc_tot_sz__10__::()>
    //***************************************************************
    //* Action task action_t3__ll_desc_tot_sz__10__
    //**************************************************************** 
   virtual task action_t3__ll_desc_tot_sz__10__(longint unsigned meta_val);
        m_t3.ll_desc_tot_sz[10] = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc_tot_sz__10__::()>

//<unsigned_meta_action::_t3__ll_desc_tot_sz__9__::()>
    //***************************************************************
    //* Action task action_t3__ll_desc_tot_sz__9__
    //**************************************************************** 
   virtual task action_t3__ll_desc_tot_sz__9__(longint unsigned meta_val);
        m_t3.ll_desc_tot_sz[9] = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc_tot_sz__9__::()>

//<unsigned_meta_action::_t3__ll_desc_tot_sz__8__::()>
    //***************************************************************
    //* Action task action_t3__ll_desc_tot_sz__8__
    //**************************************************************** 
   virtual task action_t3__ll_desc_tot_sz__8__(longint unsigned meta_val);
        m_t3.ll_desc_tot_sz[8] = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc_tot_sz__8__::()>

//<unsigned_meta_action::_t3__ll_desc_tot_sz__7__::()>
    //***************************************************************
    //* Action task action_t3__ll_desc_tot_sz__7__
    //**************************************************************** 
   virtual task action_t3__ll_desc_tot_sz__7__(longint unsigned meta_val);
        m_t3.ll_desc_tot_sz[7] = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc_tot_sz__7__::()>

//<unsigned_meta_action::_t3__ll_desc_tot_sz__6__::()>
    //***************************************************************
    //* Action task action_t3__ll_desc_tot_sz__6__
    //**************************************************************** 
   virtual task action_t3__ll_desc_tot_sz__6__(longint unsigned meta_val);
        m_t3.ll_desc_tot_sz[6] = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc_tot_sz__6__::()>

//<unsigned_meta_action::_t3__ll_desc_tot_sz__5__::()>
    //***************************************************************
    //* Action task action_t3__ll_desc_tot_sz__5__
    //**************************************************************** 
   virtual task action_t3__ll_desc_tot_sz__5__(longint unsigned meta_val);
        m_t3.ll_desc_tot_sz[5] = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc_tot_sz__5__::()>

//<unsigned_meta_action::_t3__ll_desc_tot_sz__4__::()>
    //***************************************************************
    //* Action task action_t3__ll_desc_tot_sz__4__
    //**************************************************************** 
   virtual task action_t3__ll_desc_tot_sz__4__(longint unsigned meta_val);
        m_t3.ll_desc_tot_sz[4] = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc_tot_sz__4__::()>

//<unsigned_meta_action::_t3__ll_desc_tot_sz__3__::()>
    //***************************************************************
    //* Action task action_t3__ll_desc_tot_sz__3__
    //**************************************************************** 
   virtual task action_t3__ll_desc_tot_sz__3__(longint unsigned meta_val);
        m_t3.ll_desc_tot_sz[3] = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc_tot_sz__3__::()>

//<unsigned_meta_action::_t3__ll_desc_tot_sz__2__::()>
    //***************************************************************
    //* Action task action_t3__ll_desc_tot_sz__2__
    //**************************************************************** 
   virtual task action_t3__ll_desc_tot_sz__2__(longint unsigned meta_val);
        m_t3.ll_desc_tot_sz[2] = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc_tot_sz__2__::()>

//<unsigned_meta_action::_t3__ll_desc_tot_sz__1__::()>
    //***************************************************************
    //* Action task action_t3__ll_desc_tot_sz__1__
    //**************************************************************** 
   virtual task action_t3__ll_desc_tot_sz__1__(longint unsigned meta_val);
        m_t3.ll_desc_tot_sz[1] = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc_tot_sz__1__::()>

//<unsigned_meta_action::_t3__ll_desc_tot_sz__0__::()>
    //***************************************************************
    //* Action task action_t3__ll_desc_tot_sz__0__
    //**************************************************************** 
   virtual task action_t3__ll_desc_tot_sz__0__(longint unsigned meta_val);
        m_t3.ll_desc_tot_sz[0] = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc_tot_sz__0__::()>

//<unsigned_meta_action::_t3__ll_desc_sz::()>
    //***************************************************************
    //* Action task action_t3__ll_desc_sz
    //**************************************************************** 
   virtual task action_t3__ll_desc_sz(longint unsigned meta_val);
        m_t3.ll_desc_sz = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc_sz::()>

//<unsigned_meta_action::_t3__ll_desc__15____tot_sz::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__15____tot_sz
    //**************************************************************** 
   virtual task action_t3__ll_desc__15____tot_sz(longint unsigned meta_val);
        m_t3.ll_desc[15].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__15____tot_sz::()>

//<unsigned_meta_action::_t3__ll_desc__15____dst_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__15____dst_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__15____dst_sel(longint unsigned meta_val);
        m_t3.ll_desc[15].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__15____dst_sel::()>

//<unsigned_meta_action::_t3__ll_desc__15____src_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__15____src_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__15____src_sel(longint unsigned meta_val);
        m_t3.ll_desc[15].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__15____src_sel::()>

//<unsigned_meta_action::_t3__ll_desc__15____inc_dst::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__15____inc_dst
    //**************************************************************** 
   virtual task action_t3__ll_desc__15____inc_dst(longint unsigned meta_val);
        m_t3.ll_desc[15].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__15____inc_dst::()>

//<unsigned_meta_action::_t3__ll_desc__15____inc_src::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__15____inc_src
    //**************************************************************** 
   virtual task action_t3__ll_desc__15____inc_src(longint unsigned meta_val);
        m_t3.ll_desc[15].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__15____inc_src::()>

//<unsigned_meta_action::_t3__ll_desc__14____tot_sz::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__14____tot_sz
    //**************************************************************** 
   virtual task action_t3__ll_desc__14____tot_sz(longint unsigned meta_val);
        m_t3.ll_desc[14].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__14____tot_sz::()>

//<unsigned_meta_action::_t3__ll_desc__14____dst_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__14____dst_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__14____dst_sel(longint unsigned meta_val);
        m_t3.ll_desc[14].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__14____dst_sel::()>

//<unsigned_meta_action::_t3__ll_desc__14____src_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__14____src_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__14____src_sel(longint unsigned meta_val);
        m_t3.ll_desc[14].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__14____src_sel::()>

//<unsigned_meta_action::_t3__ll_desc__14____inc_dst::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__14____inc_dst
    //**************************************************************** 
   virtual task action_t3__ll_desc__14____inc_dst(longint unsigned meta_val);
        m_t3.ll_desc[14].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__14____inc_dst::()>

//<unsigned_meta_action::_t3__ll_desc__14____inc_src::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__14____inc_src
    //**************************************************************** 
   virtual task action_t3__ll_desc__14____inc_src(longint unsigned meta_val);
        m_t3.ll_desc[14].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__14____inc_src::()>

//<unsigned_meta_action::_t3__ll_desc__13____tot_sz::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__13____tot_sz
    //**************************************************************** 
   virtual task action_t3__ll_desc__13____tot_sz(longint unsigned meta_val);
        m_t3.ll_desc[13].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__13____tot_sz::()>

//<unsigned_meta_action::_t3__ll_desc__13____dst_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__13____dst_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__13____dst_sel(longint unsigned meta_val);
        m_t3.ll_desc[13].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__13____dst_sel::()>

//<unsigned_meta_action::_t3__ll_desc__13____src_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__13____src_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__13____src_sel(longint unsigned meta_val);
        m_t3.ll_desc[13].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__13____src_sel::()>

//<unsigned_meta_action::_t3__ll_desc__13____inc_dst::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__13____inc_dst
    //**************************************************************** 
   virtual task action_t3__ll_desc__13____inc_dst(longint unsigned meta_val);
        m_t3.ll_desc[13].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__13____inc_dst::()>

//<unsigned_meta_action::_t3__ll_desc__13____inc_src::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__13____inc_src
    //**************************************************************** 
   virtual task action_t3__ll_desc__13____inc_src(longint unsigned meta_val);
        m_t3.ll_desc[13].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__13____inc_src::()>

//<unsigned_meta_action::_t3__ll_desc__12____tot_sz::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__12____tot_sz
    //**************************************************************** 
   virtual task action_t3__ll_desc__12____tot_sz(longint unsigned meta_val);
        m_t3.ll_desc[12].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__12____tot_sz::()>

//<unsigned_meta_action::_t3__ll_desc__12____dst_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__12____dst_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__12____dst_sel(longint unsigned meta_val);
        m_t3.ll_desc[12].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__12____dst_sel::()>

//<unsigned_meta_action::_t3__ll_desc__12____src_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__12____src_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__12____src_sel(longint unsigned meta_val);
        m_t3.ll_desc[12].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__12____src_sel::()>

//<unsigned_meta_action::_t3__ll_desc__12____inc_dst::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__12____inc_dst
    //**************************************************************** 
   virtual task action_t3__ll_desc__12____inc_dst(longint unsigned meta_val);
        m_t3.ll_desc[12].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__12____inc_dst::()>

//<unsigned_meta_action::_t3__ll_desc__12____inc_src::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__12____inc_src
    //**************************************************************** 
   virtual task action_t3__ll_desc__12____inc_src(longint unsigned meta_val);
        m_t3.ll_desc[12].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__12____inc_src::()>

//<unsigned_meta_action::_t3__ll_desc__11____tot_sz::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__11____tot_sz
    //**************************************************************** 
   virtual task action_t3__ll_desc__11____tot_sz(longint unsigned meta_val);
        m_t3.ll_desc[11].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__11____tot_sz::()>

//<unsigned_meta_action::_t3__ll_desc__11____dst_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__11____dst_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__11____dst_sel(longint unsigned meta_val);
        m_t3.ll_desc[11].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__11____dst_sel::()>

//<unsigned_meta_action::_t3__ll_desc__11____src_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__11____src_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__11____src_sel(longint unsigned meta_val);
        m_t3.ll_desc[11].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__11____src_sel::()>

//<unsigned_meta_action::_t3__ll_desc__11____inc_dst::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__11____inc_dst
    //**************************************************************** 
   virtual task action_t3__ll_desc__11____inc_dst(longint unsigned meta_val);
        m_t3.ll_desc[11].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__11____inc_dst::()>

//<unsigned_meta_action::_t3__ll_desc__11____inc_src::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__11____inc_src
    //**************************************************************** 
   virtual task action_t3__ll_desc__11____inc_src(longint unsigned meta_val);
        m_t3.ll_desc[11].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__11____inc_src::()>

//<unsigned_meta_action::_t3__ll_desc__10____tot_sz::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__10____tot_sz
    //**************************************************************** 
   virtual task action_t3__ll_desc__10____tot_sz(longint unsigned meta_val);
        m_t3.ll_desc[10].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__10____tot_sz::()>

//<unsigned_meta_action::_t3__ll_desc__10____dst_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__10____dst_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__10____dst_sel(longint unsigned meta_val);
        m_t3.ll_desc[10].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__10____dst_sel::()>

//<unsigned_meta_action::_t3__ll_desc__10____src_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__10____src_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__10____src_sel(longint unsigned meta_val);
        m_t3.ll_desc[10].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__10____src_sel::()>

//<unsigned_meta_action::_t3__ll_desc__10____inc_dst::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__10____inc_dst
    //**************************************************************** 
   virtual task action_t3__ll_desc__10____inc_dst(longint unsigned meta_val);
        m_t3.ll_desc[10].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__10____inc_dst::()>

//<unsigned_meta_action::_t3__ll_desc__10____inc_src::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__10____inc_src
    //**************************************************************** 
   virtual task action_t3__ll_desc__10____inc_src(longint unsigned meta_val);
        m_t3.ll_desc[10].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__10____inc_src::()>

//<unsigned_meta_action::_t3__ll_desc__9____tot_sz::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__9____tot_sz
    //**************************************************************** 
   virtual task action_t3__ll_desc__9____tot_sz(longint unsigned meta_val);
        m_t3.ll_desc[9].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__9____tot_sz::()>

//<unsigned_meta_action::_t3__ll_desc__9____dst_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__9____dst_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__9____dst_sel(longint unsigned meta_val);
        m_t3.ll_desc[9].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__9____dst_sel::()>

//<unsigned_meta_action::_t3__ll_desc__9____src_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__9____src_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__9____src_sel(longint unsigned meta_val);
        m_t3.ll_desc[9].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__9____src_sel::()>

//<unsigned_meta_action::_t3__ll_desc__9____inc_dst::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__9____inc_dst
    //**************************************************************** 
   virtual task action_t3__ll_desc__9____inc_dst(longint unsigned meta_val);
        m_t3.ll_desc[9].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__9____inc_dst::()>

//<unsigned_meta_action::_t3__ll_desc__9____inc_src::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__9____inc_src
    //**************************************************************** 
   virtual task action_t3__ll_desc__9____inc_src(longint unsigned meta_val);
        m_t3.ll_desc[9].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__9____inc_src::()>

//<unsigned_meta_action::_t3__ll_desc__8____tot_sz::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__8____tot_sz
    //**************************************************************** 
   virtual task action_t3__ll_desc__8____tot_sz(longint unsigned meta_val);
        m_t3.ll_desc[8].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__8____tot_sz::()>

//<unsigned_meta_action::_t3__ll_desc__8____dst_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__8____dst_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__8____dst_sel(longint unsigned meta_val);
        m_t3.ll_desc[8].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__8____dst_sel::()>

//<unsigned_meta_action::_t3__ll_desc__8____src_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__8____src_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__8____src_sel(longint unsigned meta_val);
        m_t3.ll_desc[8].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__8____src_sel::()>

//<unsigned_meta_action::_t3__ll_desc__8____inc_dst::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__8____inc_dst
    //**************************************************************** 
   virtual task action_t3__ll_desc__8____inc_dst(longint unsigned meta_val);
        m_t3.ll_desc[8].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__8____inc_dst::()>

//<unsigned_meta_action::_t3__ll_desc__8____inc_src::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__8____inc_src
    //**************************************************************** 
   virtual task action_t3__ll_desc__8____inc_src(longint unsigned meta_val);
        m_t3.ll_desc[8].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__8____inc_src::()>

//<unsigned_meta_action::_t3__ll_desc__7____tot_sz::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__7____tot_sz
    //**************************************************************** 
   virtual task action_t3__ll_desc__7____tot_sz(longint unsigned meta_val);
        m_t3.ll_desc[7].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__7____tot_sz::()>

//<unsigned_meta_action::_t3__ll_desc__7____dst_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__7____dst_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__7____dst_sel(longint unsigned meta_val);
        m_t3.ll_desc[7].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__7____dst_sel::()>

//<unsigned_meta_action::_t3__ll_desc__7____src_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__7____src_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__7____src_sel(longint unsigned meta_val);
        m_t3.ll_desc[7].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__7____src_sel::()>

//<unsigned_meta_action::_t3__ll_desc__7____inc_dst::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__7____inc_dst
    //**************************************************************** 
   virtual task action_t3__ll_desc__7____inc_dst(longint unsigned meta_val);
        m_t3.ll_desc[7].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__7____inc_dst::()>

//<unsigned_meta_action::_t3__ll_desc__7____inc_src::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__7____inc_src
    //**************************************************************** 
   virtual task action_t3__ll_desc__7____inc_src(longint unsigned meta_val);
        m_t3.ll_desc[7].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__7____inc_src::()>

//<unsigned_meta_action::_t3__ll_desc__6____tot_sz::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__6____tot_sz
    //**************************************************************** 
   virtual task action_t3__ll_desc__6____tot_sz(longint unsigned meta_val);
        m_t3.ll_desc[6].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__6____tot_sz::()>

//<unsigned_meta_action::_t3__ll_desc__6____dst_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__6____dst_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__6____dst_sel(longint unsigned meta_val);
        m_t3.ll_desc[6].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__6____dst_sel::()>

//<unsigned_meta_action::_t3__ll_desc__6____src_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__6____src_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__6____src_sel(longint unsigned meta_val);
        m_t3.ll_desc[6].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__6____src_sel::()>

//<unsigned_meta_action::_t3__ll_desc__6____inc_dst::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__6____inc_dst
    //**************************************************************** 
   virtual task action_t3__ll_desc__6____inc_dst(longint unsigned meta_val);
        m_t3.ll_desc[6].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__6____inc_dst::()>

//<unsigned_meta_action::_t3__ll_desc__6____inc_src::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__6____inc_src
    //**************************************************************** 
   virtual task action_t3__ll_desc__6____inc_src(longint unsigned meta_val);
        m_t3.ll_desc[6].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__6____inc_src::()>

//<unsigned_meta_action::_t3__ll_desc__5____tot_sz::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__5____tot_sz
    //**************************************************************** 
   virtual task action_t3__ll_desc__5____tot_sz(longint unsigned meta_val);
        m_t3.ll_desc[5].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__5____tot_sz::()>

//<unsigned_meta_action::_t3__ll_desc__5____dst_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__5____dst_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__5____dst_sel(longint unsigned meta_val);
        m_t3.ll_desc[5].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__5____dst_sel::()>

//<unsigned_meta_action::_t3__ll_desc__5____src_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__5____src_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__5____src_sel(longint unsigned meta_val);
        m_t3.ll_desc[5].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__5____src_sel::()>

//<unsigned_meta_action::_t3__ll_desc__5____inc_dst::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__5____inc_dst
    //**************************************************************** 
   virtual task action_t3__ll_desc__5____inc_dst(longint unsigned meta_val);
        m_t3.ll_desc[5].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__5____inc_dst::()>

//<unsigned_meta_action::_t3__ll_desc__5____inc_src::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__5____inc_src
    //**************************************************************** 
   virtual task action_t3__ll_desc__5____inc_src(longint unsigned meta_val);
        m_t3.ll_desc[5].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__5____inc_src::()>

//<unsigned_meta_action::_t3__ll_desc__4____tot_sz::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__4____tot_sz
    //**************************************************************** 
   virtual task action_t3__ll_desc__4____tot_sz(longint unsigned meta_val);
        m_t3.ll_desc[4].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__4____tot_sz::()>

//<unsigned_meta_action::_t3__ll_desc__4____dst_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__4____dst_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__4____dst_sel(longint unsigned meta_val);
        m_t3.ll_desc[4].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__4____dst_sel::()>

//<unsigned_meta_action::_t3__ll_desc__4____src_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__4____src_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__4____src_sel(longint unsigned meta_val);
        m_t3.ll_desc[4].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__4____src_sel::()>

//<unsigned_meta_action::_t3__ll_desc__4____inc_dst::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__4____inc_dst
    //**************************************************************** 
   virtual task action_t3__ll_desc__4____inc_dst(longint unsigned meta_val);
        m_t3.ll_desc[4].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__4____inc_dst::()>

//<unsigned_meta_action::_t3__ll_desc__4____inc_src::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__4____inc_src
    //**************************************************************** 
   virtual task action_t3__ll_desc__4____inc_src(longint unsigned meta_val);
        m_t3.ll_desc[4].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__4____inc_src::()>

//<unsigned_meta_action::_t3__ll_desc__3____tot_sz::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__3____tot_sz
    //**************************************************************** 
   virtual task action_t3__ll_desc__3____tot_sz(longint unsigned meta_val);
        m_t3.ll_desc[3].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__3____tot_sz::()>

//<unsigned_meta_action::_t3__ll_desc__3____dst_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__3____dst_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__3____dst_sel(longint unsigned meta_val);
        m_t3.ll_desc[3].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__3____dst_sel::()>

//<unsigned_meta_action::_t3__ll_desc__3____src_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__3____src_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__3____src_sel(longint unsigned meta_val);
        m_t3.ll_desc[3].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__3____src_sel::()>

//<unsigned_meta_action::_t3__ll_desc__3____inc_dst::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__3____inc_dst
    //**************************************************************** 
   virtual task action_t3__ll_desc__3____inc_dst(longint unsigned meta_val);
        m_t3.ll_desc[3].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__3____inc_dst::()>

//<unsigned_meta_action::_t3__ll_desc__3____inc_src::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__3____inc_src
    //**************************************************************** 
   virtual task action_t3__ll_desc__3____inc_src(longint unsigned meta_val);
        m_t3.ll_desc[3].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__3____inc_src::()>

//<unsigned_meta_action::_t3__ll_desc__2____tot_sz::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__2____tot_sz
    //**************************************************************** 
   virtual task action_t3__ll_desc__2____tot_sz(longint unsigned meta_val);
        m_t3.ll_desc[2].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__2____tot_sz::()>

//<unsigned_meta_action::_t3__ll_desc__2____dst_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__2____dst_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__2____dst_sel(longint unsigned meta_val);
        m_t3.ll_desc[2].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__2____dst_sel::()>

//<unsigned_meta_action::_t3__ll_desc__2____src_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__2____src_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__2____src_sel(longint unsigned meta_val);
        m_t3.ll_desc[2].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__2____src_sel::()>

//<unsigned_meta_action::_t3__ll_desc__2____inc_dst::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__2____inc_dst
    //**************************************************************** 
   virtual task action_t3__ll_desc__2____inc_dst(longint unsigned meta_val);
        m_t3.ll_desc[2].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__2____inc_dst::()>

//<unsigned_meta_action::_t3__ll_desc__2____inc_src::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__2____inc_src
    //**************************************************************** 
   virtual task action_t3__ll_desc__2____inc_src(longint unsigned meta_val);
        m_t3.ll_desc[2].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__2____inc_src::()>

//<unsigned_meta_action::_t3__ll_desc__1____tot_sz::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__1____tot_sz
    //**************************************************************** 
   virtual task action_t3__ll_desc__1____tot_sz(longint unsigned meta_val);
        m_t3.ll_desc[1].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__1____tot_sz::()>

//<unsigned_meta_action::_t3__ll_desc__1____dst_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__1____dst_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__1____dst_sel(longint unsigned meta_val);
        m_t3.ll_desc[1].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__1____dst_sel::()>

//<unsigned_meta_action::_t3__ll_desc__1____src_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__1____src_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__1____src_sel(longint unsigned meta_val);
        m_t3.ll_desc[1].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__1____src_sel::()>

//<unsigned_meta_action::_t3__ll_desc__1____inc_dst::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__1____inc_dst
    //**************************************************************** 
   virtual task action_t3__ll_desc__1____inc_dst(longint unsigned meta_val);
        m_t3.ll_desc[1].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__1____inc_dst::()>

//<unsigned_meta_action::_t3__ll_desc__1____inc_src::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__1____inc_src
    //**************************************************************** 
   virtual task action_t3__ll_desc__1____inc_src(longint unsigned meta_val);
        m_t3.ll_desc[1].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__1____inc_src::()>

//<unsigned_meta_action::_t3__ll_desc__0____tot_sz::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__0____tot_sz
    //**************************************************************** 
   virtual task action_t3__ll_desc__0____tot_sz(longint unsigned meta_val);
        m_t3.ll_desc[0].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__0____tot_sz::()>

//<unsigned_meta_action::_t3__ll_desc__0____dst_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__0____dst_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__0____dst_sel(longint unsigned meta_val);
        m_t3.ll_desc[0].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__0____dst_sel::()>

//<unsigned_meta_action::_t3__ll_desc__0____src_sel::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__0____src_sel
    //**************************************************************** 
   virtual task action_t3__ll_desc__0____src_sel(longint unsigned meta_val);
        m_t3.ll_desc[0].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__0____src_sel::()>

//<unsigned_meta_action::_t3__ll_desc__0____inc_dst::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__0____inc_dst
    //**************************************************************** 
   virtual task action_t3__ll_desc__0____inc_dst(longint unsigned meta_val);
        m_t3.ll_desc[0].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__0____inc_dst::()>

//<unsigned_meta_action::_t3__ll_desc__0____inc_src::()>
    //***************************************************************
    //* Action task action_t3__ll_desc__0____inc_src
    //**************************************************************** 
   virtual task action_t3__ll_desc__0____inc_src(longint unsigned meta_val);
        m_t3.ll_desc[0].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t3__ll_desc__0____inc_src::()>

//<unsigned_meta_action::_t3__chk_sz::()>
    //***************************************************************
    //* Action task action_t3__chk_sz
    //**************************************************************** 
   virtual task action_t3__chk_sz(longint unsigned meta_val);
        m_t3.chk_sz = meta_val;
    endtask
//</unsigned_meta_action::_t3__chk_sz::()>

//<unsigned_meta_action::_t3__tot_sz::()>
    //***************************************************************
    //* Action task action_t3__tot_sz
    //**************************************************************** 
   virtual task action_t3__tot_sz(longint unsigned meta_val);
        m_t3.tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t3__tot_sz::()>

//<unsigned_meta_action::_t3__dst_sel::()>
    //***************************************************************
    //* Action task action_t3__dst_sel
    //**************************************************************** 
   virtual task action_t3__dst_sel(longint unsigned meta_val);
        m_t3.dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__dst_sel::()>

//<unsigned_meta_action::_t3__src_sel::()>
    //***************************************************************
    //* Action task action_t3__src_sel
    //**************************************************************** 
   virtual task action_t3__src_sel(longint unsigned meta_val);
        m_t3.src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t3__src_sel::()>

//<unsigned_meta_action::_t3__inc_dst::()>
    //***************************************************************
    //* Action task action_t3__inc_dst
    //**************************************************************** 
   virtual task action_t3__inc_dst(longint unsigned meta_val);
        m_t3.inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t3__inc_dst::()>

//<unsigned_meta_action::_t3__inc_src::()>
    //***************************************************************
    //* Action task action_t3__inc_src
    //**************************************************************** 
   virtual task action_t3__inc_src(longint unsigned meta_val);
        m_t3.inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t3__inc_src::()>

//<unsigned_meta_action::_t3__mode::()>
    //***************************************************************
    //* Action task action_t3__mode
    //**************************************************************** 
   virtual task action_t3__mode(longint unsigned meta_val);
        m_t3.mode = meta_val;
    endtask
//</unsigned_meta_action::_t3__mode::()>

//<unsigned_meta_action::_t3__channel::()>
    //***************************************************************
    //* Action task action_t3__channel
    //**************************************************************** 
   virtual task action_t3__channel(longint unsigned meta_val);
        m_t3.channel = meta_val;
    endtask
//</unsigned_meta_action::_t3__channel::()>

//<unsigned_meta_action::_t2__transfer_sz::()>
    //***************************************************************
    //* Action task action_t2__transfer_sz
    //**************************************************************** 
   virtual task action_t2__transfer_sz(longint unsigned meta_val);
        m_t2.transfer_sz = meta_val;
    endtask
//</unsigned_meta_action::_t2__transfer_sz::()>

//<unsigned_meta_action::_t2__ll_desc_tot_sz__15__::()>
    //***************************************************************
    //* Action task action_t2__ll_desc_tot_sz__15__
    //**************************************************************** 
   virtual task action_t2__ll_desc_tot_sz__15__(longint unsigned meta_val);
        m_t2.ll_desc_tot_sz[15] = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc_tot_sz__15__::()>

//<unsigned_meta_action::_t2__ll_desc_tot_sz__14__::()>
    //***************************************************************
    //* Action task action_t2__ll_desc_tot_sz__14__
    //**************************************************************** 
   virtual task action_t2__ll_desc_tot_sz__14__(longint unsigned meta_val);
        m_t2.ll_desc_tot_sz[14] = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc_tot_sz__14__::()>

//<unsigned_meta_action::_t2__ll_desc_tot_sz__13__::()>
    //***************************************************************
    //* Action task action_t2__ll_desc_tot_sz__13__
    //**************************************************************** 
   virtual task action_t2__ll_desc_tot_sz__13__(longint unsigned meta_val);
        m_t2.ll_desc_tot_sz[13] = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc_tot_sz__13__::()>

//<unsigned_meta_action::_t2__ll_desc_tot_sz__12__::()>
    //***************************************************************
    //* Action task action_t2__ll_desc_tot_sz__12__
    //**************************************************************** 
   virtual task action_t2__ll_desc_tot_sz__12__(longint unsigned meta_val);
        m_t2.ll_desc_tot_sz[12] = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc_tot_sz__12__::()>

//<unsigned_meta_action::_t2__ll_desc_tot_sz__11__::()>
    //***************************************************************
    //* Action task action_t2__ll_desc_tot_sz__11__
    //**************************************************************** 
   virtual task action_t2__ll_desc_tot_sz__11__(longint unsigned meta_val);
        m_t2.ll_desc_tot_sz[11] = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc_tot_sz__11__::()>

//<unsigned_meta_action::_t2__ll_desc_tot_sz__10__::()>
    //***************************************************************
    //* Action task action_t2__ll_desc_tot_sz__10__
    //**************************************************************** 
   virtual task action_t2__ll_desc_tot_sz__10__(longint unsigned meta_val);
        m_t2.ll_desc_tot_sz[10] = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc_tot_sz__10__::()>

//<unsigned_meta_action::_t2__ll_desc_tot_sz__9__::()>
    //***************************************************************
    //* Action task action_t2__ll_desc_tot_sz__9__
    //**************************************************************** 
   virtual task action_t2__ll_desc_tot_sz__9__(longint unsigned meta_val);
        m_t2.ll_desc_tot_sz[9] = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc_tot_sz__9__::()>

//<unsigned_meta_action::_t2__ll_desc_tot_sz__8__::()>
    //***************************************************************
    //* Action task action_t2__ll_desc_tot_sz__8__
    //**************************************************************** 
   virtual task action_t2__ll_desc_tot_sz__8__(longint unsigned meta_val);
        m_t2.ll_desc_tot_sz[8] = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc_tot_sz__8__::()>

//<unsigned_meta_action::_t2__ll_desc_tot_sz__7__::()>
    //***************************************************************
    //* Action task action_t2__ll_desc_tot_sz__7__
    //**************************************************************** 
   virtual task action_t2__ll_desc_tot_sz__7__(longint unsigned meta_val);
        m_t2.ll_desc_tot_sz[7] = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc_tot_sz__7__::()>

//<unsigned_meta_action::_t2__ll_desc_tot_sz__6__::()>
    //***************************************************************
    //* Action task action_t2__ll_desc_tot_sz__6__
    //**************************************************************** 
   virtual task action_t2__ll_desc_tot_sz__6__(longint unsigned meta_val);
        m_t2.ll_desc_tot_sz[6] = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc_tot_sz__6__::()>

//<unsigned_meta_action::_t2__ll_desc_tot_sz__5__::()>
    //***************************************************************
    //* Action task action_t2__ll_desc_tot_sz__5__
    //**************************************************************** 
   virtual task action_t2__ll_desc_tot_sz__5__(longint unsigned meta_val);
        m_t2.ll_desc_tot_sz[5] = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc_tot_sz__5__::()>

//<unsigned_meta_action::_t2__ll_desc_tot_sz__4__::()>
    //***************************************************************
    //* Action task action_t2__ll_desc_tot_sz__4__
    //**************************************************************** 
   virtual task action_t2__ll_desc_tot_sz__4__(longint unsigned meta_val);
        m_t2.ll_desc_tot_sz[4] = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc_tot_sz__4__::()>

//<unsigned_meta_action::_t2__ll_desc_tot_sz__3__::()>
    //***************************************************************
    //* Action task action_t2__ll_desc_tot_sz__3__
    //**************************************************************** 
   virtual task action_t2__ll_desc_tot_sz__3__(longint unsigned meta_val);
        m_t2.ll_desc_tot_sz[3] = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc_tot_sz__3__::()>

//<unsigned_meta_action::_t2__ll_desc_tot_sz__2__::()>
    //***************************************************************
    //* Action task action_t2__ll_desc_tot_sz__2__
    //**************************************************************** 
   virtual task action_t2__ll_desc_tot_sz__2__(longint unsigned meta_val);
        m_t2.ll_desc_tot_sz[2] = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc_tot_sz__2__::()>

//<unsigned_meta_action::_t2__ll_desc_tot_sz__1__::()>
    //***************************************************************
    //* Action task action_t2__ll_desc_tot_sz__1__
    //**************************************************************** 
   virtual task action_t2__ll_desc_tot_sz__1__(longint unsigned meta_val);
        m_t2.ll_desc_tot_sz[1] = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc_tot_sz__1__::()>

//<unsigned_meta_action::_t2__ll_desc_tot_sz__0__::()>
    //***************************************************************
    //* Action task action_t2__ll_desc_tot_sz__0__
    //**************************************************************** 
   virtual task action_t2__ll_desc_tot_sz__0__(longint unsigned meta_val);
        m_t2.ll_desc_tot_sz[0] = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc_tot_sz__0__::()>

//<unsigned_meta_action::_t2__ll_desc_sz::()>
    //***************************************************************
    //* Action task action_t2__ll_desc_sz
    //**************************************************************** 
   virtual task action_t2__ll_desc_sz(longint unsigned meta_val);
        m_t2.ll_desc_sz = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc_sz::()>

//<unsigned_meta_action::_t2__ll_desc__15____tot_sz::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__15____tot_sz
    //**************************************************************** 
   virtual task action_t2__ll_desc__15____tot_sz(longint unsigned meta_val);
        m_t2.ll_desc[15].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__15____tot_sz::()>

//<unsigned_meta_action::_t2__ll_desc__15____dst_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__15____dst_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__15____dst_sel(longint unsigned meta_val);
        m_t2.ll_desc[15].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__15____dst_sel::()>

//<unsigned_meta_action::_t2__ll_desc__15____src_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__15____src_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__15____src_sel(longint unsigned meta_val);
        m_t2.ll_desc[15].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__15____src_sel::()>

//<unsigned_meta_action::_t2__ll_desc__15____inc_dst::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__15____inc_dst
    //**************************************************************** 
   virtual task action_t2__ll_desc__15____inc_dst(longint unsigned meta_val);
        m_t2.ll_desc[15].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__15____inc_dst::()>

//<unsigned_meta_action::_t2__ll_desc__15____inc_src::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__15____inc_src
    //**************************************************************** 
   virtual task action_t2__ll_desc__15____inc_src(longint unsigned meta_val);
        m_t2.ll_desc[15].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__15____inc_src::()>

//<unsigned_meta_action::_t2__ll_desc__14____tot_sz::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__14____tot_sz
    //**************************************************************** 
   virtual task action_t2__ll_desc__14____tot_sz(longint unsigned meta_val);
        m_t2.ll_desc[14].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__14____tot_sz::()>

//<unsigned_meta_action::_t2__ll_desc__14____dst_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__14____dst_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__14____dst_sel(longint unsigned meta_val);
        m_t2.ll_desc[14].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__14____dst_sel::()>

//<unsigned_meta_action::_t2__ll_desc__14____src_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__14____src_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__14____src_sel(longint unsigned meta_val);
        m_t2.ll_desc[14].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__14____src_sel::()>

//<unsigned_meta_action::_t2__ll_desc__14____inc_dst::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__14____inc_dst
    //**************************************************************** 
   virtual task action_t2__ll_desc__14____inc_dst(longint unsigned meta_val);
        m_t2.ll_desc[14].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__14____inc_dst::()>

//<unsigned_meta_action::_t2__ll_desc__14____inc_src::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__14____inc_src
    //**************************************************************** 
   virtual task action_t2__ll_desc__14____inc_src(longint unsigned meta_val);
        m_t2.ll_desc[14].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__14____inc_src::()>

//<unsigned_meta_action::_t2__ll_desc__13____tot_sz::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__13____tot_sz
    //**************************************************************** 
   virtual task action_t2__ll_desc__13____tot_sz(longint unsigned meta_val);
        m_t2.ll_desc[13].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__13____tot_sz::()>

//<unsigned_meta_action::_t2__ll_desc__13____dst_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__13____dst_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__13____dst_sel(longint unsigned meta_val);
        m_t2.ll_desc[13].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__13____dst_sel::()>

//<unsigned_meta_action::_t2__ll_desc__13____src_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__13____src_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__13____src_sel(longint unsigned meta_val);
        m_t2.ll_desc[13].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__13____src_sel::()>

//<unsigned_meta_action::_t2__ll_desc__13____inc_dst::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__13____inc_dst
    //**************************************************************** 
   virtual task action_t2__ll_desc__13____inc_dst(longint unsigned meta_val);
        m_t2.ll_desc[13].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__13____inc_dst::()>

//<unsigned_meta_action::_t2__ll_desc__13____inc_src::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__13____inc_src
    //**************************************************************** 
   virtual task action_t2__ll_desc__13____inc_src(longint unsigned meta_val);
        m_t2.ll_desc[13].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__13____inc_src::()>

//<unsigned_meta_action::_t2__ll_desc__12____tot_sz::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__12____tot_sz
    //**************************************************************** 
   virtual task action_t2__ll_desc__12____tot_sz(longint unsigned meta_val);
        m_t2.ll_desc[12].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__12____tot_sz::()>

//<unsigned_meta_action::_t2__ll_desc__12____dst_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__12____dst_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__12____dst_sel(longint unsigned meta_val);
        m_t2.ll_desc[12].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__12____dst_sel::()>

//<unsigned_meta_action::_t2__ll_desc__12____src_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__12____src_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__12____src_sel(longint unsigned meta_val);
        m_t2.ll_desc[12].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__12____src_sel::()>

//<unsigned_meta_action::_t2__ll_desc__12____inc_dst::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__12____inc_dst
    //**************************************************************** 
   virtual task action_t2__ll_desc__12____inc_dst(longint unsigned meta_val);
        m_t2.ll_desc[12].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__12____inc_dst::()>

//<unsigned_meta_action::_t2__ll_desc__12____inc_src::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__12____inc_src
    //**************************************************************** 
   virtual task action_t2__ll_desc__12____inc_src(longint unsigned meta_val);
        m_t2.ll_desc[12].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__12____inc_src::()>

//<unsigned_meta_action::_t2__ll_desc__11____tot_sz::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__11____tot_sz
    //**************************************************************** 
   virtual task action_t2__ll_desc__11____tot_sz(longint unsigned meta_val);
        m_t2.ll_desc[11].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__11____tot_sz::()>

//<unsigned_meta_action::_t2__ll_desc__11____dst_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__11____dst_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__11____dst_sel(longint unsigned meta_val);
        m_t2.ll_desc[11].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__11____dst_sel::()>

//<unsigned_meta_action::_t2__ll_desc__11____src_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__11____src_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__11____src_sel(longint unsigned meta_val);
        m_t2.ll_desc[11].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__11____src_sel::()>

//<unsigned_meta_action::_t2__ll_desc__11____inc_dst::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__11____inc_dst
    //**************************************************************** 
   virtual task action_t2__ll_desc__11____inc_dst(longint unsigned meta_val);
        m_t2.ll_desc[11].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__11____inc_dst::()>

//<unsigned_meta_action::_t2__ll_desc__11____inc_src::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__11____inc_src
    //**************************************************************** 
   virtual task action_t2__ll_desc__11____inc_src(longint unsigned meta_val);
        m_t2.ll_desc[11].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__11____inc_src::()>

//<unsigned_meta_action::_t2__ll_desc__10____tot_sz::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__10____tot_sz
    //**************************************************************** 
   virtual task action_t2__ll_desc__10____tot_sz(longint unsigned meta_val);
        m_t2.ll_desc[10].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__10____tot_sz::()>

//<unsigned_meta_action::_t2__ll_desc__10____dst_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__10____dst_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__10____dst_sel(longint unsigned meta_val);
        m_t2.ll_desc[10].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__10____dst_sel::()>

//<unsigned_meta_action::_t2__ll_desc__10____src_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__10____src_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__10____src_sel(longint unsigned meta_val);
        m_t2.ll_desc[10].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__10____src_sel::()>

//<unsigned_meta_action::_t2__ll_desc__10____inc_dst::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__10____inc_dst
    //**************************************************************** 
   virtual task action_t2__ll_desc__10____inc_dst(longint unsigned meta_val);
        m_t2.ll_desc[10].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__10____inc_dst::()>

//<unsigned_meta_action::_t2__ll_desc__10____inc_src::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__10____inc_src
    //**************************************************************** 
   virtual task action_t2__ll_desc__10____inc_src(longint unsigned meta_val);
        m_t2.ll_desc[10].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__10____inc_src::()>

//<unsigned_meta_action::_t2__ll_desc__9____tot_sz::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__9____tot_sz
    //**************************************************************** 
   virtual task action_t2__ll_desc__9____tot_sz(longint unsigned meta_val);
        m_t2.ll_desc[9].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__9____tot_sz::()>

//<unsigned_meta_action::_t2__ll_desc__9____dst_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__9____dst_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__9____dst_sel(longint unsigned meta_val);
        m_t2.ll_desc[9].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__9____dst_sel::()>

//<unsigned_meta_action::_t2__ll_desc__9____src_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__9____src_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__9____src_sel(longint unsigned meta_val);
        m_t2.ll_desc[9].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__9____src_sel::()>

//<unsigned_meta_action::_t2__ll_desc__9____inc_dst::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__9____inc_dst
    //**************************************************************** 
   virtual task action_t2__ll_desc__9____inc_dst(longint unsigned meta_val);
        m_t2.ll_desc[9].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__9____inc_dst::()>

//<unsigned_meta_action::_t2__ll_desc__9____inc_src::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__9____inc_src
    //**************************************************************** 
   virtual task action_t2__ll_desc__9____inc_src(longint unsigned meta_val);
        m_t2.ll_desc[9].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__9____inc_src::()>

//<unsigned_meta_action::_t2__ll_desc__8____tot_sz::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__8____tot_sz
    //**************************************************************** 
   virtual task action_t2__ll_desc__8____tot_sz(longint unsigned meta_val);
        m_t2.ll_desc[8].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__8____tot_sz::()>

//<unsigned_meta_action::_t2__ll_desc__8____dst_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__8____dst_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__8____dst_sel(longint unsigned meta_val);
        m_t2.ll_desc[8].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__8____dst_sel::()>

//<unsigned_meta_action::_t2__ll_desc__8____src_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__8____src_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__8____src_sel(longint unsigned meta_val);
        m_t2.ll_desc[8].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__8____src_sel::()>

//<unsigned_meta_action::_t2__ll_desc__8____inc_dst::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__8____inc_dst
    //**************************************************************** 
   virtual task action_t2__ll_desc__8____inc_dst(longint unsigned meta_val);
        m_t2.ll_desc[8].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__8____inc_dst::()>

//<unsigned_meta_action::_t2__ll_desc__8____inc_src::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__8____inc_src
    //**************************************************************** 
   virtual task action_t2__ll_desc__8____inc_src(longint unsigned meta_val);
        m_t2.ll_desc[8].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__8____inc_src::()>

//<unsigned_meta_action::_t2__ll_desc__7____tot_sz::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__7____tot_sz
    //**************************************************************** 
   virtual task action_t2__ll_desc__7____tot_sz(longint unsigned meta_val);
        m_t2.ll_desc[7].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__7____tot_sz::()>

//<unsigned_meta_action::_t2__ll_desc__7____dst_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__7____dst_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__7____dst_sel(longint unsigned meta_val);
        m_t2.ll_desc[7].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__7____dst_sel::()>

//<unsigned_meta_action::_t2__ll_desc__7____src_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__7____src_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__7____src_sel(longint unsigned meta_val);
        m_t2.ll_desc[7].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__7____src_sel::()>

//<unsigned_meta_action::_t2__ll_desc__7____inc_dst::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__7____inc_dst
    //**************************************************************** 
   virtual task action_t2__ll_desc__7____inc_dst(longint unsigned meta_val);
        m_t2.ll_desc[7].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__7____inc_dst::()>

//<unsigned_meta_action::_t2__ll_desc__7____inc_src::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__7____inc_src
    //**************************************************************** 
   virtual task action_t2__ll_desc__7____inc_src(longint unsigned meta_val);
        m_t2.ll_desc[7].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__7____inc_src::()>

//<unsigned_meta_action::_t2__ll_desc__6____tot_sz::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__6____tot_sz
    //**************************************************************** 
   virtual task action_t2__ll_desc__6____tot_sz(longint unsigned meta_val);
        m_t2.ll_desc[6].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__6____tot_sz::()>

//<unsigned_meta_action::_t2__ll_desc__6____dst_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__6____dst_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__6____dst_sel(longint unsigned meta_val);
        m_t2.ll_desc[6].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__6____dst_sel::()>

//<unsigned_meta_action::_t2__ll_desc__6____src_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__6____src_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__6____src_sel(longint unsigned meta_val);
        m_t2.ll_desc[6].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__6____src_sel::()>

//<unsigned_meta_action::_t2__ll_desc__6____inc_dst::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__6____inc_dst
    //**************************************************************** 
   virtual task action_t2__ll_desc__6____inc_dst(longint unsigned meta_val);
        m_t2.ll_desc[6].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__6____inc_dst::()>

//<unsigned_meta_action::_t2__ll_desc__6____inc_src::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__6____inc_src
    //**************************************************************** 
   virtual task action_t2__ll_desc__6____inc_src(longint unsigned meta_val);
        m_t2.ll_desc[6].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__6____inc_src::()>

//<unsigned_meta_action::_t2__ll_desc__5____tot_sz::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__5____tot_sz
    //**************************************************************** 
   virtual task action_t2__ll_desc__5____tot_sz(longint unsigned meta_val);
        m_t2.ll_desc[5].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__5____tot_sz::()>

//<unsigned_meta_action::_t2__ll_desc__5____dst_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__5____dst_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__5____dst_sel(longint unsigned meta_val);
        m_t2.ll_desc[5].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__5____dst_sel::()>

//<unsigned_meta_action::_t2__ll_desc__5____src_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__5____src_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__5____src_sel(longint unsigned meta_val);
        m_t2.ll_desc[5].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__5____src_sel::()>

//<unsigned_meta_action::_t2__ll_desc__5____inc_dst::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__5____inc_dst
    //**************************************************************** 
   virtual task action_t2__ll_desc__5____inc_dst(longint unsigned meta_val);
        m_t2.ll_desc[5].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__5____inc_dst::()>

//<unsigned_meta_action::_t2__ll_desc__5____inc_src::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__5____inc_src
    //**************************************************************** 
   virtual task action_t2__ll_desc__5____inc_src(longint unsigned meta_val);
        m_t2.ll_desc[5].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__5____inc_src::()>

//<unsigned_meta_action::_t2__ll_desc__4____tot_sz::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__4____tot_sz
    //**************************************************************** 
   virtual task action_t2__ll_desc__4____tot_sz(longint unsigned meta_val);
        m_t2.ll_desc[4].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__4____tot_sz::()>

//<unsigned_meta_action::_t2__ll_desc__4____dst_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__4____dst_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__4____dst_sel(longint unsigned meta_val);
        m_t2.ll_desc[4].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__4____dst_sel::()>

//<unsigned_meta_action::_t2__ll_desc__4____src_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__4____src_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__4____src_sel(longint unsigned meta_val);
        m_t2.ll_desc[4].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__4____src_sel::()>

//<unsigned_meta_action::_t2__ll_desc__4____inc_dst::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__4____inc_dst
    //**************************************************************** 
   virtual task action_t2__ll_desc__4____inc_dst(longint unsigned meta_val);
        m_t2.ll_desc[4].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__4____inc_dst::()>

//<unsigned_meta_action::_t2__ll_desc__4____inc_src::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__4____inc_src
    //**************************************************************** 
   virtual task action_t2__ll_desc__4____inc_src(longint unsigned meta_val);
        m_t2.ll_desc[4].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__4____inc_src::()>

//<unsigned_meta_action::_t2__ll_desc__3____tot_sz::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__3____tot_sz
    //**************************************************************** 
   virtual task action_t2__ll_desc__3____tot_sz(longint unsigned meta_val);
        m_t2.ll_desc[3].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__3____tot_sz::()>

//<unsigned_meta_action::_t2__ll_desc__3____dst_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__3____dst_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__3____dst_sel(longint unsigned meta_val);
        m_t2.ll_desc[3].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__3____dst_sel::()>

//<unsigned_meta_action::_t2__ll_desc__3____src_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__3____src_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__3____src_sel(longint unsigned meta_val);
        m_t2.ll_desc[3].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__3____src_sel::()>

//<unsigned_meta_action::_t2__ll_desc__3____inc_dst::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__3____inc_dst
    //**************************************************************** 
   virtual task action_t2__ll_desc__3____inc_dst(longint unsigned meta_val);
        m_t2.ll_desc[3].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__3____inc_dst::()>

//<unsigned_meta_action::_t2__ll_desc__3____inc_src::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__3____inc_src
    //**************************************************************** 
   virtual task action_t2__ll_desc__3____inc_src(longint unsigned meta_val);
        m_t2.ll_desc[3].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__3____inc_src::()>

//<unsigned_meta_action::_t2__ll_desc__2____tot_sz::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__2____tot_sz
    //**************************************************************** 
   virtual task action_t2__ll_desc__2____tot_sz(longint unsigned meta_val);
        m_t2.ll_desc[2].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__2____tot_sz::()>

//<unsigned_meta_action::_t2__ll_desc__2____dst_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__2____dst_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__2____dst_sel(longint unsigned meta_val);
        m_t2.ll_desc[2].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__2____dst_sel::()>

//<unsigned_meta_action::_t2__ll_desc__2____src_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__2____src_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__2____src_sel(longint unsigned meta_val);
        m_t2.ll_desc[2].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__2____src_sel::()>

//<unsigned_meta_action::_t2__ll_desc__2____inc_dst::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__2____inc_dst
    //**************************************************************** 
   virtual task action_t2__ll_desc__2____inc_dst(longint unsigned meta_val);
        m_t2.ll_desc[2].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__2____inc_dst::()>

//<unsigned_meta_action::_t2__ll_desc__2____inc_src::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__2____inc_src
    //**************************************************************** 
   virtual task action_t2__ll_desc__2____inc_src(longint unsigned meta_val);
        m_t2.ll_desc[2].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__2____inc_src::()>

//<unsigned_meta_action::_t2__ll_desc__1____tot_sz::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__1____tot_sz
    //**************************************************************** 
   virtual task action_t2__ll_desc__1____tot_sz(longint unsigned meta_val);
        m_t2.ll_desc[1].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__1____tot_sz::()>

//<unsigned_meta_action::_t2__ll_desc__1____dst_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__1____dst_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__1____dst_sel(longint unsigned meta_val);
        m_t2.ll_desc[1].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__1____dst_sel::()>

//<unsigned_meta_action::_t2__ll_desc__1____src_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__1____src_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__1____src_sel(longint unsigned meta_val);
        m_t2.ll_desc[1].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__1____src_sel::()>

//<unsigned_meta_action::_t2__ll_desc__1____inc_dst::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__1____inc_dst
    //**************************************************************** 
   virtual task action_t2__ll_desc__1____inc_dst(longint unsigned meta_val);
        m_t2.ll_desc[1].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__1____inc_dst::()>

//<unsigned_meta_action::_t2__ll_desc__1____inc_src::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__1____inc_src
    //**************************************************************** 
   virtual task action_t2__ll_desc__1____inc_src(longint unsigned meta_val);
        m_t2.ll_desc[1].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__1____inc_src::()>

//<unsigned_meta_action::_t2__ll_desc__0____tot_sz::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__0____tot_sz
    //**************************************************************** 
   virtual task action_t2__ll_desc__0____tot_sz(longint unsigned meta_val);
        m_t2.ll_desc[0].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__0____tot_sz::()>

//<unsigned_meta_action::_t2__ll_desc__0____dst_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__0____dst_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__0____dst_sel(longint unsigned meta_val);
        m_t2.ll_desc[0].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__0____dst_sel::()>

//<unsigned_meta_action::_t2__ll_desc__0____src_sel::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__0____src_sel
    //**************************************************************** 
   virtual task action_t2__ll_desc__0____src_sel(longint unsigned meta_val);
        m_t2.ll_desc[0].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__0____src_sel::()>

//<unsigned_meta_action::_t2__ll_desc__0____inc_dst::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__0____inc_dst
    //**************************************************************** 
   virtual task action_t2__ll_desc__0____inc_dst(longint unsigned meta_val);
        m_t2.ll_desc[0].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__0____inc_dst::()>

//<unsigned_meta_action::_t2__ll_desc__0____inc_src::()>
    //***************************************************************
    //* Action task action_t2__ll_desc__0____inc_src
    //**************************************************************** 
   virtual task action_t2__ll_desc__0____inc_src(longint unsigned meta_val);
        m_t2.ll_desc[0].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t2__ll_desc__0____inc_src::()>

//<unsigned_meta_action::_t2__chk_sz::()>
    //***************************************************************
    //* Action task action_t2__chk_sz
    //**************************************************************** 
   virtual task action_t2__chk_sz(longint unsigned meta_val);
        m_t2.chk_sz = meta_val;
    endtask
//</unsigned_meta_action::_t2__chk_sz::()>

//<unsigned_meta_action::_t2__tot_sz::()>
    //***************************************************************
    //* Action task action_t2__tot_sz
    //**************************************************************** 
   virtual task action_t2__tot_sz(longint unsigned meta_val);
        m_t2.tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t2__tot_sz::()>

//<unsigned_meta_action::_t2__dst_sel::()>
    //***************************************************************
    //* Action task action_t2__dst_sel
    //**************************************************************** 
   virtual task action_t2__dst_sel(longint unsigned meta_val);
        m_t2.dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__dst_sel::()>

//<unsigned_meta_action::_t2__src_sel::()>
    //***************************************************************
    //* Action task action_t2__src_sel
    //**************************************************************** 
   virtual task action_t2__src_sel(longint unsigned meta_val);
        m_t2.src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t2__src_sel::()>

//<unsigned_meta_action::_t2__inc_dst::()>
    //***************************************************************
    //* Action task action_t2__inc_dst
    //**************************************************************** 
   virtual task action_t2__inc_dst(longint unsigned meta_val);
        m_t2.inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t2__inc_dst::()>

//<unsigned_meta_action::_t2__inc_src::()>
    //***************************************************************
    //* Action task action_t2__inc_src
    //**************************************************************** 
   virtual task action_t2__inc_src(longint unsigned meta_val);
        m_t2.inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t2__inc_src::()>

//<unsigned_meta_action::_t2__mode::()>
    //***************************************************************
    //* Action task action_t2__mode
    //**************************************************************** 
   virtual task action_t2__mode(longint unsigned meta_val);
        m_t2.mode = meta_val;
    endtask
//</unsigned_meta_action::_t2__mode::()>

//<unsigned_meta_action::_t2__channel::()>
    //***************************************************************
    //* Action task action_t2__channel
    //**************************************************************** 
   virtual task action_t2__channel(longint unsigned meta_val);
        m_t2.channel = meta_val;
    endtask
//</unsigned_meta_action::_t2__channel::()>

//<unsigned_meta_action::_t1__transfer_sz::()>
    //***************************************************************
    //* Action task action_t1__transfer_sz
    //**************************************************************** 
   virtual task action_t1__transfer_sz(longint unsigned meta_val);
        m_t1.transfer_sz = meta_val;
    endtask
//</unsigned_meta_action::_t1__transfer_sz::()>

//<unsigned_meta_action::_t1__ll_desc_tot_sz__15__::()>
    //***************************************************************
    //* Action task action_t1__ll_desc_tot_sz__15__
    //**************************************************************** 
   virtual task action_t1__ll_desc_tot_sz__15__(longint unsigned meta_val);
        m_t1.ll_desc_tot_sz[15] = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc_tot_sz__15__::()>

//<unsigned_meta_action::_t1__ll_desc_tot_sz__14__::()>
    //***************************************************************
    //* Action task action_t1__ll_desc_tot_sz__14__
    //**************************************************************** 
   virtual task action_t1__ll_desc_tot_sz__14__(longint unsigned meta_val);
        m_t1.ll_desc_tot_sz[14] = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc_tot_sz__14__::()>

//<unsigned_meta_action::_t1__ll_desc_tot_sz__13__::()>
    //***************************************************************
    //* Action task action_t1__ll_desc_tot_sz__13__
    //**************************************************************** 
   virtual task action_t1__ll_desc_tot_sz__13__(longint unsigned meta_val);
        m_t1.ll_desc_tot_sz[13] = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc_tot_sz__13__::()>

//<unsigned_meta_action::_t1__ll_desc_tot_sz__12__::()>
    //***************************************************************
    //* Action task action_t1__ll_desc_tot_sz__12__
    //**************************************************************** 
   virtual task action_t1__ll_desc_tot_sz__12__(longint unsigned meta_val);
        m_t1.ll_desc_tot_sz[12] = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc_tot_sz__12__::()>

//<unsigned_meta_action::_t1__ll_desc_tot_sz__11__::()>
    //***************************************************************
    //* Action task action_t1__ll_desc_tot_sz__11__
    //**************************************************************** 
   virtual task action_t1__ll_desc_tot_sz__11__(longint unsigned meta_val);
        m_t1.ll_desc_tot_sz[11] = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc_tot_sz__11__::()>

//<unsigned_meta_action::_t1__ll_desc_tot_sz__10__::()>
    //***************************************************************
    //* Action task action_t1__ll_desc_tot_sz__10__
    //**************************************************************** 
   virtual task action_t1__ll_desc_tot_sz__10__(longint unsigned meta_val);
        m_t1.ll_desc_tot_sz[10] = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc_tot_sz__10__::()>

//<unsigned_meta_action::_t1__ll_desc_tot_sz__9__::()>
    //***************************************************************
    //* Action task action_t1__ll_desc_tot_sz__9__
    //**************************************************************** 
   virtual task action_t1__ll_desc_tot_sz__9__(longint unsigned meta_val);
        m_t1.ll_desc_tot_sz[9] = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc_tot_sz__9__::()>

//<unsigned_meta_action::_t1__ll_desc_tot_sz__8__::()>
    //***************************************************************
    //* Action task action_t1__ll_desc_tot_sz__8__
    //**************************************************************** 
   virtual task action_t1__ll_desc_tot_sz__8__(longint unsigned meta_val);
        m_t1.ll_desc_tot_sz[8] = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc_tot_sz__8__::()>

//<unsigned_meta_action::_t1__ll_desc_tot_sz__7__::()>
    //***************************************************************
    //* Action task action_t1__ll_desc_tot_sz__7__
    //**************************************************************** 
   virtual task action_t1__ll_desc_tot_sz__7__(longint unsigned meta_val);
        m_t1.ll_desc_tot_sz[7] = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc_tot_sz__7__::()>

//<unsigned_meta_action::_t1__ll_desc_tot_sz__6__::()>
    //***************************************************************
    //* Action task action_t1__ll_desc_tot_sz__6__
    //**************************************************************** 
   virtual task action_t1__ll_desc_tot_sz__6__(longint unsigned meta_val);
        m_t1.ll_desc_tot_sz[6] = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc_tot_sz__6__::()>

//<unsigned_meta_action::_t1__ll_desc_tot_sz__5__::()>
    //***************************************************************
    //* Action task action_t1__ll_desc_tot_sz__5__
    //**************************************************************** 
   virtual task action_t1__ll_desc_tot_sz__5__(longint unsigned meta_val);
        m_t1.ll_desc_tot_sz[5] = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc_tot_sz__5__::()>

//<unsigned_meta_action::_t1__ll_desc_tot_sz__4__::()>
    //***************************************************************
    //* Action task action_t1__ll_desc_tot_sz__4__
    //**************************************************************** 
   virtual task action_t1__ll_desc_tot_sz__4__(longint unsigned meta_val);
        m_t1.ll_desc_tot_sz[4] = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc_tot_sz__4__::()>

//<unsigned_meta_action::_t1__ll_desc_tot_sz__3__::()>
    //***************************************************************
    //* Action task action_t1__ll_desc_tot_sz__3__
    //**************************************************************** 
   virtual task action_t1__ll_desc_tot_sz__3__(longint unsigned meta_val);
        m_t1.ll_desc_tot_sz[3] = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc_tot_sz__3__::()>

//<unsigned_meta_action::_t1__ll_desc_tot_sz__2__::()>
    //***************************************************************
    //* Action task action_t1__ll_desc_tot_sz__2__
    //**************************************************************** 
   virtual task action_t1__ll_desc_tot_sz__2__(longint unsigned meta_val);
        m_t1.ll_desc_tot_sz[2] = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc_tot_sz__2__::()>

//<unsigned_meta_action::_t1__ll_desc_tot_sz__1__::()>
    //***************************************************************
    //* Action task action_t1__ll_desc_tot_sz__1__
    //**************************************************************** 
   virtual task action_t1__ll_desc_tot_sz__1__(longint unsigned meta_val);
        m_t1.ll_desc_tot_sz[1] = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc_tot_sz__1__::()>

//<unsigned_meta_action::_t1__ll_desc_tot_sz__0__::()>
    //***************************************************************
    //* Action task action_t1__ll_desc_tot_sz__0__
    //**************************************************************** 
   virtual task action_t1__ll_desc_tot_sz__0__(longint unsigned meta_val);
        m_t1.ll_desc_tot_sz[0] = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc_tot_sz__0__::()>

//<unsigned_meta_action::_t1__ll_desc_sz::()>
    //***************************************************************
    //* Action task action_t1__ll_desc_sz
    //**************************************************************** 
   virtual task action_t1__ll_desc_sz(longint unsigned meta_val);
        m_t1.ll_desc_sz = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc_sz::()>

//<unsigned_meta_action::_t1__ll_desc__15____tot_sz::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__15____tot_sz
    //**************************************************************** 
   virtual task action_t1__ll_desc__15____tot_sz(longint unsigned meta_val);
        m_t1.ll_desc[15].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__15____tot_sz::()>

//<unsigned_meta_action::_t1__ll_desc__15____dst_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__15____dst_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__15____dst_sel(longint unsigned meta_val);
        m_t1.ll_desc[15].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__15____dst_sel::()>

//<unsigned_meta_action::_t1__ll_desc__15____src_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__15____src_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__15____src_sel(longint unsigned meta_val);
        m_t1.ll_desc[15].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__15____src_sel::()>

//<unsigned_meta_action::_t1__ll_desc__15____inc_dst::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__15____inc_dst
    //**************************************************************** 
   virtual task action_t1__ll_desc__15____inc_dst(longint unsigned meta_val);
        m_t1.ll_desc[15].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__15____inc_dst::()>

//<unsigned_meta_action::_t1__ll_desc__15____inc_src::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__15____inc_src
    //**************************************************************** 
   virtual task action_t1__ll_desc__15____inc_src(longint unsigned meta_val);
        m_t1.ll_desc[15].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__15____inc_src::()>

//<unsigned_meta_action::_t1__ll_desc__14____tot_sz::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__14____tot_sz
    //**************************************************************** 
   virtual task action_t1__ll_desc__14____tot_sz(longint unsigned meta_val);
        m_t1.ll_desc[14].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__14____tot_sz::()>

//<unsigned_meta_action::_t1__ll_desc__14____dst_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__14____dst_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__14____dst_sel(longint unsigned meta_val);
        m_t1.ll_desc[14].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__14____dst_sel::()>

//<unsigned_meta_action::_t1__ll_desc__14____src_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__14____src_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__14____src_sel(longint unsigned meta_val);
        m_t1.ll_desc[14].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__14____src_sel::()>

//<unsigned_meta_action::_t1__ll_desc__14____inc_dst::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__14____inc_dst
    //**************************************************************** 
   virtual task action_t1__ll_desc__14____inc_dst(longint unsigned meta_val);
        m_t1.ll_desc[14].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__14____inc_dst::()>

//<unsigned_meta_action::_t1__ll_desc__14____inc_src::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__14____inc_src
    //**************************************************************** 
   virtual task action_t1__ll_desc__14____inc_src(longint unsigned meta_val);
        m_t1.ll_desc[14].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__14____inc_src::()>

//<unsigned_meta_action::_t1__ll_desc__13____tot_sz::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__13____tot_sz
    //**************************************************************** 
   virtual task action_t1__ll_desc__13____tot_sz(longint unsigned meta_val);
        m_t1.ll_desc[13].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__13____tot_sz::()>

//<unsigned_meta_action::_t1__ll_desc__13____dst_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__13____dst_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__13____dst_sel(longint unsigned meta_val);
        m_t1.ll_desc[13].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__13____dst_sel::()>

//<unsigned_meta_action::_t1__ll_desc__13____src_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__13____src_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__13____src_sel(longint unsigned meta_val);
        m_t1.ll_desc[13].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__13____src_sel::()>

//<unsigned_meta_action::_t1__ll_desc__13____inc_dst::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__13____inc_dst
    //**************************************************************** 
   virtual task action_t1__ll_desc__13____inc_dst(longint unsigned meta_val);
        m_t1.ll_desc[13].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__13____inc_dst::()>

//<unsigned_meta_action::_t1__ll_desc__13____inc_src::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__13____inc_src
    //**************************************************************** 
   virtual task action_t1__ll_desc__13____inc_src(longint unsigned meta_val);
        m_t1.ll_desc[13].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__13____inc_src::()>

//<unsigned_meta_action::_t1__ll_desc__12____tot_sz::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__12____tot_sz
    //**************************************************************** 
   virtual task action_t1__ll_desc__12____tot_sz(longint unsigned meta_val);
        m_t1.ll_desc[12].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__12____tot_sz::()>

//<unsigned_meta_action::_t1__ll_desc__12____dst_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__12____dst_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__12____dst_sel(longint unsigned meta_val);
        m_t1.ll_desc[12].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__12____dst_sel::()>

//<unsigned_meta_action::_t1__ll_desc__12____src_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__12____src_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__12____src_sel(longint unsigned meta_val);
        m_t1.ll_desc[12].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__12____src_sel::()>

//<unsigned_meta_action::_t1__ll_desc__12____inc_dst::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__12____inc_dst
    //**************************************************************** 
   virtual task action_t1__ll_desc__12____inc_dst(longint unsigned meta_val);
        m_t1.ll_desc[12].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__12____inc_dst::()>

//<unsigned_meta_action::_t1__ll_desc__12____inc_src::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__12____inc_src
    //**************************************************************** 
   virtual task action_t1__ll_desc__12____inc_src(longint unsigned meta_val);
        m_t1.ll_desc[12].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__12____inc_src::()>

//<unsigned_meta_action::_t1__ll_desc__11____tot_sz::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__11____tot_sz
    //**************************************************************** 
   virtual task action_t1__ll_desc__11____tot_sz(longint unsigned meta_val);
        m_t1.ll_desc[11].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__11____tot_sz::()>

//<unsigned_meta_action::_t1__ll_desc__11____dst_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__11____dst_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__11____dst_sel(longint unsigned meta_val);
        m_t1.ll_desc[11].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__11____dst_sel::()>

//<unsigned_meta_action::_t1__ll_desc__11____src_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__11____src_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__11____src_sel(longint unsigned meta_val);
        m_t1.ll_desc[11].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__11____src_sel::()>

//<unsigned_meta_action::_t1__ll_desc__11____inc_dst::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__11____inc_dst
    //**************************************************************** 
   virtual task action_t1__ll_desc__11____inc_dst(longint unsigned meta_val);
        m_t1.ll_desc[11].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__11____inc_dst::()>

//<unsigned_meta_action::_t1__ll_desc__11____inc_src::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__11____inc_src
    //**************************************************************** 
   virtual task action_t1__ll_desc__11____inc_src(longint unsigned meta_val);
        m_t1.ll_desc[11].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__11____inc_src::()>

//<unsigned_meta_action::_t1__ll_desc__10____tot_sz::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__10____tot_sz
    //**************************************************************** 
   virtual task action_t1__ll_desc__10____tot_sz(longint unsigned meta_val);
        m_t1.ll_desc[10].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__10____tot_sz::()>

//<unsigned_meta_action::_t1__ll_desc__10____dst_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__10____dst_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__10____dst_sel(longint unsigned meta_val);
        m_t1.ll_desc[10].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__10____dst_sel::()>

//<unsigned_meta_action::_t1__ll_desc__10____src_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__10____src_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__10____src_sel(longint unsigned meta_val);
        m_t1.ll_desc[10].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__10____src_sel::()>

//<unsigned_meta_action::_t1__ll_desc__10____inc_dst::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__10____inc_dst
    //**************************************************************** 
   virtual task action_t1__ll_desc__10____inc_dst(longint unsigned meta_val);
        m_t1.ll_desc[10].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__10____inc_dst::()>

//<unsigned_meta_action::_t1__ll_desc__10____inc_src::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__10____inc_src
    //**************************************************************** 
   virtual task action_t1__ll_desc__10____inc_src(longint unsigned meta_val);
        m_t1.ll_desc[10].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__10____inc_src::()>

//<unsigned_meta_action::_t1__ll_desc__9____tot_sz::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__9____tot_sz
    //**************************************************************** 
   virtual task action_t1__ll_desc__9____tot_sz(longint unsigned meta_val);
        m_t1.ll_desc[9].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__9____tot_sz::()>

//<unsigned_meta_action::_t1__ll_desc__9____dst_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__9____dst_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__9____dst_sel(longint unsigned meta_val);
        m_t1.ll_desc[9].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__9____dst_sel::()>

//<unsigned_meta_action::_t1__ll_desc__9____src_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__9____src_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__9____src_sel(longint unsigned meta_val);
        m_t1.ll_desc[9].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__9____src_sel::()>

//<unsigned_meta_action::_t1__ll_desc__9____inc_dst::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__9____inc_dst
    //**************************************************************** 
   virtual task action_t1__ll_desc__9____inc_dst(longint unsigned meta_val);
        m_t1.ll_desc[9].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__9____inc_dst::()>

//<unsigned_meta_action::_t1__ll_desc__9____inc_src::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__9____inc_src
    //**************************************************************** 
   virtual task action_t1__ll_desc__9____inc_src(longint unsigned meta_val);
        m_t1.ll_desc[9].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__9____inc_src::()>

//<unsigned_meta_action::_t1__ll_desc__8____tot_sz::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__8____tot_sz
    //**************************************************************** 
   virtual task action_t1__ll_desc__8____tot_sz(longint unsigned meta_val);
        m_t1.ll_desc[8].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__8____tot_sz::()>

//<unsigned_meta_action::_t1__ll_desc__8____dst_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__8____dst_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__8____dst_sel(longint unsigned meta_val);
        m_t1.ll_desc[8].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__8____dst_sel::()>

//<unsigned_meta_action::_t1__ll_desc__8____src_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__8____src_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__8____src_sel(longint unsigned meta_val);
        m_t1.ll_desc[8].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__8____src_sel::()>

//<unsigned_meta_action::_t1__ll_desc__8____inc_dst::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__8____inc_dst
    //**************************************************************** 
   virtual task action_t1__ll_desc__8____inc_dst(longint unsigned meta_val);
        m_t1.ll_desc[8].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__8____inc_dst::()>

//<unsigned_meta_action::_t1__ll_desc__8____inc_src::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__8____inc_src
    //**************************************************************** 
   virtual task action_t1__ll_desc__8____inc_src(longint unsigned meta_val);
        m_t1.ll_desc[8].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__8____inc_src::()>

//<unsigned_meta_action::_t1__ll_desc__7____tot_sz::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__7____tot_sz
    //**************************************************************** 
   virtual task action_t1__ll_desc__7____tot_sz(longint unsigned meta_val);
        m_t1.ll_desc[7].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__7____tot_sz::()>

//<unsigned_meta_action::_t1__ll_desc__7____dst_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__7____dst_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__7____dst_sel(longint unsigned meta_val);
        m_t1.ll_desc[7].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__7____dst_sel::()>

//<unsigned_meta_action::_t1__ll_desc__7____src_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__7____src_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__7____src_sel(longint unsigned meta_val);
        m_t1.ll_desc[7].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__7____src_sel::()>

//<unsigned_meta_action::_t1__ll_desc__7____inc_dst::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__7____inc_dst
    //**************************************************************** 
   virtual task action_t1__ll_desc__7____inc_dst(longint unsigned meta_val);
        m_t1.ll_desc[7].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__7____inc_dst::()>

//<unsigned_meta_action::_t1__ll_desc__7____inc_src::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__7____inc_src
    //**************************************************************** 
   virtual task action_t1__ll_desc__7____inc_src(longint unsigned meta_val);
        m_t1.ll_desc[7].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__7____inc_src::()>

//<unsigned_meta_action::_t1__ll_desc__6____tot_sz::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__6____tot_sz
    //**************************************************************** 
   virtual task action_t1__ll_desc__6____tot_sz(longint unsigned meta_val);
        m_t1.ll_desc[6].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__6____tot_sz::()>

//<unsigned_meta_action::_t1__ll_desc__6____dst_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__6____dst_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__6____dst_sel(longint unsigned meta_val);
        m_t1.ll_desc[6].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__6____dst_sel::()>

//<unsigned_meta_action::_t1__ll_desc__6____src_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__6____src_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__6____src_sel(longint unsigned meta_val);
        m_t1.ll_desc[6].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__6____src_sel::()>

//<unsigned_meta_action::_t1__ll_desc__6____inc_dst::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__6____inc_dst
    //**************************************************************** 
   virtual task action_t1__ll_desc__6____inc_dst(longint unsigned meta_val);
        m_t1.ll_desc[6].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__6____inc_dst::()>

//<unsigned_meta_action::_t1__ll_desc__6____inc_src::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__6____inc_src
    //**************************************************************** 
   virtual task action_t1__ll_desc__6____inc_src(longint unsigned meta_val);
        m_t1.ll_desc[6].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__6____inc_src::()>

//<unsigned_meta_action::_t1__ll_desc__5____tot_sz::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__5____tot_sz
    //**************************************************************** 
   virtual task action_t1__ll_desc__5____tot_sz(longint unsigned meta_val);
        m_t1.ll_desc[5].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__5____tot_sz::()>

//<unsigned_meta_action::_t1__ll_desc__5____dst_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__5____dst_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__5____dst_sel(longint unsigned meta_val);
        m_t1.ll_desc[5].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__5____dst_sel::()>

//<unsigned_meta_action::_t1__ll_desc__5____src_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__5____src_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__5____src_sel(longint unsigned meta_val);
        m_t1.ll_desc[5].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__5____src_sel::()>

//<unsigned_meta_action::_t1__ll_desc__5____inc_dst::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__5____inc_dst
    //**************************************************************** 
   virtual task action_t1__ll_desc__5____inc_dst(longint unsigned meta_val);
        m_t1.ll_desc[5].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__5____inc_dst::()>

//<unsigned_meta_action::_t1__ll_desc__5____inc_src::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__5____inc_src
    //**************************************************************** 
   virtual task action_t1__ll_desc__5____inc_src(longint unsigned meta_val);
        m_t1.ll_desc[5].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__5____inc_src::()>

//<unsigned_meta_action::_t1__ll_desc__4____tot_sz::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__4____tot_sz
    //**************************************************************** 
   virtual task action_t1__ll_desc__4____tot_sz(longint unsigned meta_val);
        m_t1.ll_desc[4].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__4____tot_sz::()>

//<unsigned_meta_action::_t1__ll_desc__4____dst_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__4____dst_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__4____dst_sel(longint unsigned meta_val);
        m_t1.ll_desc[4].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__4____dst_sel::()>

//<unsigned_meta_action::_t1__ll_desc__4____src_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__4____src_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__4____src_sel(longint unsigned meta_val);
        m_t1.ll_desc[4].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__4____src_sel::()>

//<unsigned_meta_action::_t1__ll_desc__4____inc_dst::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__4____inc_dst
    //**************************************************************** 
   virtual task action_t1__ll_desc__4____inc_dst(longint unsigned meta_val);
        m_t1.ll_desc[4].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__4____inc_dst::()>

//<unsigned_meta_action::_t1__ll_desc__4____inc_src::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__4____inc_src
    //**************************************************************** 
   virtual task action_t1__ll_desc__4____inc_src(longint unsigned meta_val);
        m_t1.ll_desc[4].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__4____inc_src::()>

//<unsigned_meta_action::_t1__ll_desc__3____tot_sz::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__3____tot_sz
    //**************************************************************** 
   virtual task action_t1__ll_desc__3____tot_sz(longint unsigned meta_val);
        m_t1.ll_desc[3].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__3____tot_sz::()>

//<unsigned_meta_action::_t1__ll_desc__3____dst_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__3____dst_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__3____dst_sel(longint unsigned meta_val);
        m_t1.ll_desc[3].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__3____dst_sel::()>

//<unsigned_meta_action::_t1__ll_desc__3____src_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__3____src_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__3____src_sel(longint unsigned meta_val);
        m_t1.ll_desc[3].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__3____src_sel::()>

//<unsigned_meta_action::_t1__ll_desc__3____inc_dst::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__3____inc_dst
    //**************************************************************** 
   virtual task action_t1__ll_desc__3____inc_dst(longint unsigned meta_val);
        m_t1.ll_desc[3].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__3____inc_dst::()>

//<unsigned_meta_action::_t1__ll_desc__3____inc_src::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__3____inc_src
    //**************************************************************** 
   virtual task action_t1__ll_desc__3____inc_src(longint unsigned meta_val);
        m_t1.ll_desc[3].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__3____inc_src::()>

//<unsigned_meta_action::_t1__ll_desc__2____tot_sz::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__2____tot_sz
    //**************************************************************** 
   virtual task action_t1__ll_desc__2____tot_sz(longint unsigned meta_val);
        m_t1.ll_desc[2].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__2____tot_sz::()>

//<unsigned_meta_action::_t1__ll_desc__2____dst_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__2____dst_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__2____dst_sel(longint unsigned meta_val);
        m_t1.ll_desc[2].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__2____dst_sel::()>

//<unsigned_meta_action::_t1__ll_desc__2____src_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__2____src_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__2____src_sel(longint unsigned meta_val);
        m_t1.ll_desc[2].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__2____src_sel::()>

//<unsigned_meta_action::_t1__ll_desc__2____inc_dst::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__2____inc_dst
    //**************************************************************** 
   virtual task action_t1__ll_desc__2____inc_dst(longint unsigned meta_val);
        m_t1.ll_desc[2].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__2____inc_dst::()>

//<unsigned_meta_action::_t1__ll_desc__2____inc_src::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__2____inc_src
    //**************************************************************** 
   virtual task action_t1__ll_desc__2____inc_src(longint unsigned meta_val);
        m_t1.ll_desc[2].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__2____inc_src::()>

//<unsigned_meta_action::_t1__ll_desc__1____tot_sz::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__1____tot_sz
    //**************************************************************** 
   virtual task action_t1__ll_desc__1____tot_sz(longint unsigned meta_val);
        m_t1.ll_desc[1].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__1____tot_sz::()>

//<unsigned_meta_action::_t1__ll_desc__1____dst_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__1____dst_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__1____dst_sel(longint unsigned meta_val);
        m_t1.ll_desc[1].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__1____dst_sel::()>

//<unsigned_meta_action::_t1__ll_desc__1____src_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__1____src_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__1____src_sel(longint unsigned meta_val);
        m_t1.ll_desc[1].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__1____src_sel::()>

//<unsigned_meta_action::_t1__ll_desc__1____inc_dst::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__1____inc_dst
    //**************************************************************** 
   virtual task action_t1__ll_desc__1____inc_dst(longint unsigned meta_val);
        m_t1.ll_desc[1].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__1____inc_dst::()>

//<unsigned_meta_action::_t1__ll_desc__1____inc_src::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__1____inc_src
    //**************************************************************** 
   virtual task action_t1__ll_desc__1____inc_src(longint unsigned meta_val);
        m_t1.ll_desc[1].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__1____inc_src::()>

//<unsigned_meta_action::_t1__ll_desc__0____tot_sz::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__0____tot_sz
    //**************************************************************** 
   virtual task action_t1__ll_desc__0____tot_sz(longint unsigned meta_val);
        m_t1.ll_desc[0].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__0____tot_sz::()>

//<unsigned_meta_action::_t1__ll_desc__0____dst_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__0____dst_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__0____dst_sel(longint unsigned meta_val);
        m_t1.ll_desc[0].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__0____dst_sel::()>

//<unsigned_meta_action::_t1__ll_desc__0____src_sel::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__0____src_sel
    //**************************************************************** 
   virtual task action_t1__ll_desc__0____src_sel(longint unsigned meta_val);
        m_t1.ll_desc[0].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__0____src_sel::()>

//<unsigned_meta_action::_t1__ll_desc__0____inc_dst::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__0____inc_dst
    //**************************************************************** 
   virtual task action_t1__ll_desc__0____inc_dst(longint unsigned meta_val);
        m_t1.ll_desc[0].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__0____inc_dst::()>

//<unsigned_meta_action::_t1__ll_desc__0____inc_src::()>
    //***************************************************************
    //* Action task action_t1__ll_desc__0____inc_src
    //**************************************************************** 
   virtual task action_t1__ll_desc__0____inc_src(longint unsigned meta_val);
        m_t1.ll_desc[0].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t1__ll_desc__0____inc_src::()>

//<unsigned_meta_action::_t1__chk_sz::()>
    //***************************************************************
    //* Action task action_t1__chk_sz
    //**************************************************************** 
   virtual task action_t1__chk_sz(longint unsigned meta_val);
        m_t1.chk_sz = meta_val;
    endtask
//</unsigned_meta_action::_t1__chk_sz::()>

//<unsigned_meta_action::_t1__tot_sz::()>
    //***************************************************************
    //* Action task action_t1__tot_sz
    //**************************************************************** 
   virtual task action_t1__tot_sz(longint unsigned meta_val);
        m_t1.tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_t1__tot_sz::()>

//<unsigned_meta_action::_t1__dst_sel::()>
    //***************************************************************
    //* Action task action_t1__dst_sel
    //**************************************************************** 
   virtual task action_t1__dst_sel(longint unsigned meta_val);
        m_t1.dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__dst_sel::()>

//<unsigned_meta_action::_t1__src_sel::()>
    //***************************************************************
    //* Action task action_t1__src_sel
    //**************************************************************** 
   virtual task action_t1__src_sel(longint unsigned meta_val);
        m_t1.src_sel = meta_val;
    endtask
//</unsigned_meta_action::_t1__src_sel::()>

//<unsigned_meta_action::_t1__inc_dst::()>
    //***************************************************************
    //* Action task action_t1__inc_dst
    //**************************************************************** 
   virtual task action_t1__inc_dst(longint unsigned meta_val);
        m_t1.inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_t1__inc_dst::()>

//<unsigned_meta_action::_t1__inc_src::()>
    //***************************************************************
    //* Action task action_t1__inc_src
    //**************************************************************** 
   virtual task action_t1__inc_src(longint unsigned meta_val);
        m_t1.inc_src = meta_val;
    endtask
//</unsigned_meta_action::_t1__inc_src::()>

//<unsigned_meta_action::_t1__mode::()>
    //***************************************************************
    //* Action task action_t1__mode
    //**************************************************************** 
   virtual task action_t1__mode(longint unsigned meta_val);
        m_t1.mode = meta_val;
    endtask
//</unsigned_meta_action::_t1__mode::()>

//<unsigned_meta_action::_t1__channel::()>
    //***************************************************************
    //* Action task action_t1__channel
    //**************************************************************** 
   virtual task action_t1__channel(longint unsigned meta_val);
        m_t1.channel = meta_val;
    endtask
//</unsigned_meta_action::_t1__channel::()>

//<action::_wait_done::(##58bded9f0416a01b395ff75ecdd9b2c0)>
    //***************************************************************
    //* Action task action_wait_done
    //* action_stmt = wait_done();
    //**************************************************************** 
   virtual task action_wait_done();
        wait_done();
    endtask
//</action::_wait_done::(##58bded9f0416a01b395ff75ecdd9b2c0)>

//</action_tasks>
    
//<cov_cb_functions>
    /****************************************************************
     * Coverage Callback Functions
     ****************************************************************/

	/****************************************************************
	 * pathCoverageCallback() 
	 ****************************************************************/
	function void pathCoverageCallback(PathCoverage pc, CoverageCallbackReason reason);
		if (reason == Covered) begin
			$display("Path Coverage %s Complete", pc.name());
		end
	endfunction
//</cov_cb_functions>

//<end_of_replay>
	virtual function void end_of_replay();
	  m_replayEndReached = 1;
	endfunction
//</end_of_replay>

//<cov_create_functions>

//<create_cov_strategies,gen>
    function void create_cov_strategies();
    m_pc_closure = new(this);


    endfunction
//</create_cov_strategies>

//<coverage_check_report_methods,gen>
   	function string getCoverageReport();
		string report = "";
		
		return report;
	endfunction
		
	function bit allCoverageGoalsHaveBeenMet();
		bit met = 1;
		int n_checked = 0;

		return (met && n_checked > 0);
	endfunction    	
//</coverage_check_report_methods>

//</cov_create_functions>
    
    /****************************************************************
     * Private Class Methods
     ****************************************************************/
//<graph_extern,gen>
	extern function int get_graph_trace_option(string instance_name);
//</graph_extern>

     
    /**
     * register_actions()
     *
     * Register action tasks with the scheduler 
     *
     */     
    extern function void register_actions();

endclass

// Implementation of the register_actions function
`include "wb_dma_infact_4par_sw_seq_register_actions.svh"

`endif /* INCLUDED_wb_dma_infact_4par_sw_seq_SVH */

`ifdef UNDEFINED
//<trashcan,gen>
//<action::_do_item__wb_dma_infact_4par_sw_seq_item_c_inst__end::()>
    //***************************************************************
    //* Action task action_do_item__wb_dma_infact_4par_sw_seq_item_c_inst__end
    //**************************************************************** 
   virtual task action_do_item__wb_dma_infact_4par_sw_seq_item_c_inst__end();
                if (m_terminateOnReplayEnd && m_replayEndReached) begin
          `uvm_info(get_full_name(), "Skipping finish_item due to replay end", UVM_MEDIUM);
        end else begin
          finish_item(m_wb_dma_infact_4par_sw_seq_item_c_inst);
        end

    endtask
//</action::_do_item__wb_dma_infact_4par_sw_seq_item_c_inst__end::()>
//<action::_do_item__wb_dma_infact_4par_sw_seq_item_c_inst__begin::()>
    //***************************************************************
    //* Action task action_do_item__wb_dma_infact_4par_sw_seq_item_c_inst__begin
    //**************************************************************** 
   virtual task action_do_item__wb_dma_infact_4par_sw_seq_item_c_inst__begin();
        m_wb_dma_infact_4par_sw_seq_item_c_inst = wb_dma_infact_4par_sw_seq_item_c::type_id::create();
        if (m_terminateOnReplayEnd && m_replayEndReached) begin
          `uvm_info(get_full_name(), "Skipping start_item due to replay end", UVM_MEDIUM);
        end else begin
          start_item(m_wb_dma_infact_4par_sw_seq_item_c_inst);
        end

    endtask
//</action::_do_item__wb_dma_infact_4par_sw_seq_item_c_inst__begin::()>
//<action::_init::()>
    //***************************************************************
    //* Action task action_init
    //**************************************************************** 
   virtual task action_init();
    endtask
//</action::_init::()>
//<action::_xfer_4par__wait_done::()>
    //***************************************************************
    //* Action task action_xfer_4par__wait_done
    //**************************************************************** 
   virtual task action_xfer_4par__wait_done();
    endtask
//</action::_xfer_4par__wait_done::()>
//<action::_init_xfer__xfer_4par__t4__end::()>
    //***************************************************************
    //* Action task action_init_xfer__xfer_4par__t4__end
    //**************************************************************** 
   virtual task action_init_xfer__xfer_4par__t4__end();
                if (m_terminateOnReplayEnd && m_replayEndReached) begin
          `uvm_info(get_full_name(), "Skipping finish_item due to replay end", UVM_MEDIUM);
        end else begin
          finish_item(m_xfer_4par__t4);
        end

    endtask
//</action::_init_xfer__xfer_4par__t4__end::()>
//<action::_init_xfer__xfer_4par__t4__begin::()>
    //***************************************************************
    //* Action task action_init_xfer__xfer_4par__t4__begin
    //**************************************************************** 
   virtual task action_init_xfer__xfer_4par__t4__begin();
        m_xfer_4par__t4 = wb_dma_descriptor::type_id::create();
        if (m_terminateOnReplayEnd && m_replayEndReached) begin
          `uvm_info(get_full_name(), "Skipping start_item due to replay end", UVM_MEDIUM);
        end else begin
          start_item(m_xfer_4par__t4);
        end

    endtask
//</action::_init_xfer__xfer_4par__t4__begin::()>
//<action::_init_xfer__xfer_4par__t3__end::()>
    //***************************************************************
    //* Action task action_init_xfer__xfer_4par__t3__end
    //**************************************************************** 
   virtual task action_init_xfer__xfer_4par__t3__end();
                if (m_terminateOnReplayEnd && m_replayEndReached) begin
          `uvm_info(get_full_name(), "Skipping finish_item due to replay end", UVM_MEDIUM);
        end else begin
          finish_item(m_xfer_4par__t3);
        end

    endtask
//</action::_init_xfer__xfer_4par__t3__end::()>
//<action::_init_xfer__xfer_4par__t3__begin::()>
    //***************************************************************
    //* Action task action_init_xfer__xfer_4par__t3__begin
    //**************************************************************** 
   virtual task action_init_xfer__xfer_4par__t3__begin();
        m_xfer_4par__t3 = wb_dma_descriptor::type_id::create();
        if (m_terminateOnReplayEnd && m_replayEndReached) begin
          `uvm_info(get_full_name(), "Skipping start_item due to replay end", UVM_MEDIUM);
        end else begin
          start_item(m_xfer_4par__t3);
        end

    endtask
//</action::_init_xfer__xfer_4par__t3__begin::()>
//<action::_init_xfer__xfer_4par__t2__end::()>
    //***************************************************************
    //* Action task action_init_xfer__xfer_4par__t2__end
    //**************************************************************** 
   virtual task action_init_xfer__xfer_4par__t2__end();
                if (m_terminateOnReplayEnd && m_replayEndReached) begin
          `uvm_info(get_full_name(), "Skipping finish_item due to replay end", UVM_MEDIUM);
        end else begin
          finish_item(m_xfer_4par__t2);
        end

    endtask
//</action::_init_xfer__xfer_4par__t2__end::()>
//<action::_init_xfer__xfer_4par__t2__begin::()>
    //***************************************************************
    //* Action task action_init_xfer__xfer_4par__t2__begin
    //**************************************************************** 
   virtual task action_init_xfer__xfer_4par__t2__begin();
        m_xfer_4par__t2 = wb_dma_descriptor::type_id::create();
        if (m_terminateOnReplayEnd && m_replayEndReached) begin
          `uvm_info(get_full_name(), "Skipping start_item due to replay end", UVM_MEDIUM);
        end else begin
          start_item(m_xfer_4par__t2);
        end

    endtask
//</action::_init_xfer__xfer_4par__t2__begin::()>
//<action::_init_xfer__xfer_4par__t1__end::()>
    //***************************************************************
    //* Action task action_init_xfer__xfer_4par__t1__end
    //**************************************************************** 
   virtual task action_init_xfer__xfer_4par__t1__end();
                if (m_terminateOnReplayEnd && m_replayEndReached) begin
          `uvm_info(get_full_name(), "Skipping finish_item due to replay end", UVM_MEDIUM);
        end else begin
          finish_item(m_xfer_4par__t1);
        end

    endtask
//</action::_init_xfer__xfer_4par__t1__end::()>
//<action::_init_xfer__xfer_4par__t1__begin::()>
    //***************************************************************
    //* Action task action_init_xfer__xfer_4par__t1__begin
    //**************************************************************** 
   virtual task action_init_xfer__xfer_4par__t1__begin();
        m_xfer_4par__t1 = wb_dma_descriptor::type_id::create();
        if (m_terminateOnReplayEnd && m_replayEndReached) begin
          `uvm_info(get_full_name(), "Skipping start_item due to replay end", UVM_MEDIUM);
        end else begin
          start_item(m_xfer_4par__t1);
        end

    endtask
//</action::_init_xfer__xfer_4par__t1__begin::()>
//<signed_meta_action::_xfer_4par__t4__ll_desc_tot_sz__sum::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc_tot_sz__sum
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc_tot_sz__sum(longint meta_val);
        m_xfer_4par__t4__ll_desc_tot_sz__sum = meta_val;
    endtask
//</signed_meta_action::_xfer_4par__t4__ll_desc_tot_sz__sum::()>
//<signed_meta_action::_xfer_4par__t3__ll_desc_tot_sz__sum::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc_tot_sz__sum
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc_tot_sz__sum(longint meta_val);
        m_xfer_4par__t3__ll_desc_tot_sz__sum = meta_val;
    endtask
//</signed_meta_action::_xfer_4par__t3__ll_desc_tot_sz__sum::()>
//<signed_meta_action::_xfer_4par__t2__ll_desc_tot_sz__sum::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc_tot_sz__sum
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc_tot_sz__sum(longint meta_val);
        m_xfer_4par__t2__ll_desc_tot_sz__sum = meta_val;
    endtask
//</signed_meta_action::_xfer_4par__t2__ll_desc_tot_sz__sum::()>
//<signed_meta_action::_xfer_4par__t1__ll_desc_tot_sz__sum::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc_tot_sz__sum
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc_tot_sz__sum(longint meta_val);
        m_xfer_4par__t1__ll_desc_tot_sz__sum = meta_val;
    endtask
//</signed_meta_action::_xfer_4par__t1__ll_desc_tot_sz__sum::()>
//<unsigned_meta_action::_xfer_4par__t4__transfer_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__transfer_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t4__transfer_sz(longint unsigned meta_val);
        m_xfer_4par.t4.transfer_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__transfer_sz::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__15__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc_tot_sz__15__
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc_tot_sz__15__(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc_tot_sz[15] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__15__::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__14__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc_tot_sz__14__
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc_tot_sz__14__(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc_tot_sz[14] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__14__::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__13__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc_tot_sz__13__
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc_tot_sz__13__(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc_tot_sz[13] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__13__::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__12__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc_tot_sz__12__
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc_tot_sz__12__(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc_tot_sz[12] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__12__::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__11__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc_tot_sz__11__
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc_tot_sz__11__(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc_tot_sz[11] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__11__::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__10__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc_tot_sz__10__
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc_tot_sz__10__(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc_tot_sz[10] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__10__::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__9__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc_tot_sz__9__
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc_tot_sz__9__(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc_tot_sz[9] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__9__::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__8__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc_tot_sz__8__
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc_tot_sz__8__(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc_tot_sz[8] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__8__::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__7__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc_tot_sz__7__
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc_tot_sz__7__(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc_tot_sz[7] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__7__::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__6__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc_tot_sz__6__
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc_tot_sz__6__(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc_tot_sz[6] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__6__::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__5__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc_tot_sz__5__
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc_tot_sz__5__(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc_tot_sz[5] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__5__::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__4__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc_tot_sz__4__
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc_tot_sz__4__(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc_tot_sz[4] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__4__::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__3__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc_tot_sz__3__
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc_tot_sz__3__(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc_tot_sz[3] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__3__::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__2__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc_tot_sz__2__
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc_tot_sz__2__(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc_tot_sz[2] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__2__::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__1__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc_tot_sz__1__
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc_tot_sz__1__(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc_tot_sz[1] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__1__::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__0__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc_tot_sz__0__
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc_tot_sz__0__(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc_tot_sz[0] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc_tot_sz__0__::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc_sz(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc_sz::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__15____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__15____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__15____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[15].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__15____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__15____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__15____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__15____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[15].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__15____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__15____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__15____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__15____src_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[15].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__15____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__15____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__15____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__15____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[15].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__15____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__15____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__15____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__15____inc_src(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[15].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__15____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__14____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__14____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__14____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[14].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__14____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__14____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__14____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__14____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[14].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__14____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__14____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__14____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__14____src_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[14].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__14____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__14____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__14____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__14____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[14].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__14____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__14____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__14____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__14____inc_src(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[14].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__14____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__13____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__13____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__13____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[13].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__13____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__13____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__13____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__13____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[13].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__13____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__13____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__13____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__13____src_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[13].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__13____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__13____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__13____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__13____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[13].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__13____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__13____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__13____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__13____inc_src(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[13].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__13____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__12____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__12____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__12____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[12].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__12____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__12____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__12____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__12____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[12].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__12____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__12____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__12____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__12____src_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[12].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__12____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__12____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__12____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__12____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[12].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__12____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__12____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__12____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__12____inc_src(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[12].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__12____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__11____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__11____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__11____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[11].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__11____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__11____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__11____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__11____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[11].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__11____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__11____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__11____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__11____src_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[11].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__11____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__11____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__11____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__11____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[11].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__11____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__11____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__11____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__11____inc_src(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[11].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__11____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__10____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__10____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__10____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[10].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__10____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__10____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__10____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__10____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[10].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__10____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__10____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__10____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__10____src_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[10].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__10____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__10____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__10____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__10____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[10].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__10____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__10____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__10____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__10____inc_src(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[10].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__10____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__9____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__9____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__9____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[9].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__9____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__9____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__9____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__9____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[9].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__9____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__9____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__9____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__9____src_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[9].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__9____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__9____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__9____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__9____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[9].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__9____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__9____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__9____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__9____inc_src(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[9].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__9____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__8____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__8____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__8____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[8].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__8____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__8____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__8____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__8____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[8].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__8____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__8____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__8____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__8____src_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[8].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__8____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__8____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__8____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__8____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[8].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__8____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__8____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__8____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__8____inc_src(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[8].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__8____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__7____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__7____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__7____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[7].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__7____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__7____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__7____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__7____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[7].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__7____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__7____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__7____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__7____src_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[7].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__7____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__7____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__7____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__7____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[7].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__7____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__7____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__7____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__7____inc_src(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[7].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__7____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__6____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__6____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__6____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[6].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__6____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__6____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__6____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__6____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[6].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__6____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__6____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__6____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__6____src_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[6].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__6____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__6____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__6____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__6____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[6].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__6____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__6____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__6____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__6____inc_src(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[6].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__6____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__5____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__5____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__5____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[5].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__5____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__5____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__5____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__5____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[5].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__5____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__5____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__5____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__5____src_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[5].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__5____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__5____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__5____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__5____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[5].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__5____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__5____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__5____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__5____inc_src(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[5].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__5____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__4____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__4____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__4____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[4].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__4____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__4____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__4____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__4____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[4].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__4____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__4____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__4____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__4____src_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[4].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__4____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__4____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__4____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__4____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[4].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__4____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__4____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__4____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__4____inc_src(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[4].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__4____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__3____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__3____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__3____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[3].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__3____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__3____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__3____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__3____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[3].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__3____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__3____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__3____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__3____src_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[3].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__3____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__3____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__3____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__3____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[3].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__3____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__3____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__3____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__3____inc_src(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[3].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__3____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__2____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__2____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__2____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[2].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__2____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__2____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__2____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__2____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[2].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__2____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__2____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__2____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__2____src_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[2].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__2____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__2____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__2____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__2____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[2].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__2____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__2____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__2____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__2____inc_src(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[2].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__2____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__1____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__1____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__1____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[1].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__1____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__1____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__1____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__1____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[1].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__1____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__1____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__1____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__1____src_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[1].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__1____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__1____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__1____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__1____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[1].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__1____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__1____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__1____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__1____inc_src(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[1].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__1____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__0____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__0____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__0____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[0].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__0____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__0____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__0____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__0____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[0].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__0____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__0____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__0____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__0____src_sel(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[0].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__0____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__0____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__0____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__0____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[0].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__0____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t4__ll_desc__0____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__ll_desc__0____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t4__ll_desc__0____inc_src(longint unsigned meta_val);
        m_xfer_4par.t4.ll_desc[0].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__ll_desc__0____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t4__chk_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__chk_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t4__chk_sz(longint unsigned meta_val);
        m_xfer_4par.t4.chk_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__chk_sz::()>
//<unsigned_meta_action::_xfer_4par__t4__tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t4__tot_sz(longint unsigned meta_val);
        m_xfer_4par.t4.tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t4__dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__dst_sel(longint unsigned meta_val);
        m_xfer_4par.t4.dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__src_sel(longint unsigned meta_val);
        m_xfer_4par.t4.src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__src_sel::()>
//<unsigned_meta_action::_xfer_4par__t4__inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t4__inc_dst(longint unsigned meta_val);
        m_xfer_4par.t4.inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t4__inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t4__inc_src(longint unsigned meta_val);
        m_xfer_4par.t4.inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__inc_src::()>
//<unsigned_meta_action::_xfer_4par__t4__mode::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__mode
    //**************************************************************** 
   virtual task action_xfer_4par__t4__mode(longint unsigned meta_val);
        m_xfer_4par.t4.mode = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__mode::()>
//<unsigned_meta_action::_xfer_4par__t4__channel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t4__channel
    //**************************************************************** 
   virtual task action_xfer_4par__t4__channel(longint unsigned meta_val);
        m_xfer_4par.t4.channel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t4__channel::()>
//<unsigned_meta_action::_xfer_4par__t3__transfer_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__transfer_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t3__transfer_sz(longint unsigned meta_val);
        m_xfer_4par.t3.transfer_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__transfer_sz::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__15__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc_tot_sz__15__
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc_tot_sz__15__(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc_tot_sz[15] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__15__::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__14__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc_tot_sz__14__
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc_tot_sz__14__(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc_tot_sz[14] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__14__::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__13__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc_tot_sz__13__
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc_tot_sz__13__(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc_tot_sz[13] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__13__::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__12__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc_tot_sz__12__
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc_tot_sz__12__(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc_tot_sz[12] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__12__::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__11__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc_tot_sz__11__
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc_tot_sz__11__(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc_tot_sz[11] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__11__::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__10__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc_tot_sz__10__
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc_tot_sz__10__(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc_tot_sz[10] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__10__::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__9__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc_tot_sz__9__
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc_tot_sz__9__(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc_tot_sz[9] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__9__::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__8__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc_tot_sz__8__
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc_tot_sz__8__(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc_tot_sz[8] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__8__::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__7__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc_tot_sz__7__
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc_tot_sz__7__(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc_tot_sz[7] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__7__::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__6__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc_tot_sz__6__
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc_tot_sz__6__(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc_tot_sz[6] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__6__::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__5__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc_tot_sz__5__
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc_tot_sz__5__(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc_tot_sz[5] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__5__::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__4__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc_tot_sz__4__
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc_tot_sz__4__(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc_tot_sz[4] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__4__::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__3__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc_tot_sz__3__
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc_tot_sz__3__(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc_tot_sz[3] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__3__::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__2__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc_tot_sz__2__
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc_tot_sz__2__(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc_tot_sz[2] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__2__::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__1__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc_tot_sz__1__
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc_tot_sz__1__(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc_tot_sz[1] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__1__::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__0__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc_tot_sz__0__
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc_tot_sz__0__(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc_tot_sz[0] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc_tot_sz__0__::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc_sz(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc_sz::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__15____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__15____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__15____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[15].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__15____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__15____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__15____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__15____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[15].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__15____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__15____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__15____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__15____src_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[15].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__15____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__15____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__15____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__15____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[15].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__15____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__15____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__15____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__15____inc_src(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[15].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__15____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__14____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__14____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__14____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[14].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__14____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__14____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__14____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__14____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[14].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__14____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__14____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__14____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__14____src_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[14].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__14____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__14____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__14____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__14____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[14].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__14____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__14____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__14____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__14____inc_src(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[14].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__14____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__13____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__13____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__13____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[13].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__13____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__13____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__13____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__13____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[13].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__13____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__13____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__13____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__13____src_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[13].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__13____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__13____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__13____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__13____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[13].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__13____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__13____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__13____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__13____inc_src(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[13].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__13____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__12____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__12____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__12____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[12].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__12____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__12____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__12____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__12____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[12].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__12____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__12____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__12____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__12____src_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[12].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__12____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__12____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__12____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__12____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[12].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__12____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__12____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__12____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__12____inc_src(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[12].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__12____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__11____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__11____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__11____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[11].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__11____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__11____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__11____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__11____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[11].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__11____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__11____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__11____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__11____src_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[11].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__11____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__11____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__11____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__11____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[11].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__11____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__11____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__11____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__11____inc_src(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[11].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__11____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__10____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__10____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__10____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[10].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__10____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__10____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__10____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__10____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[10].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__10____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__10____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__10____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__10____src_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[10].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__10____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__10____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__10____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__10____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[10].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__10____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__10____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__10____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__10____inc_src(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[10].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__10____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__9____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__9____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__9____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[9].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__9____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__9____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__9____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__9____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[9].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__9____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__9____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__9____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__9____src_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[9].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__9____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__9____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__9____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__9____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[9].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__9____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__9____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__9____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__9____inc_src(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[9].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__9____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__8____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__8____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__8____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[8].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__8____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__8____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__8____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__8____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[8].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__8____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__8____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__8____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__8____src_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[8].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__8____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__8____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__8____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__8____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[8].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__8____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__8____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__8____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__8____inc_src(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[8].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__8____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__7____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__7____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__7____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[7].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__7____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__7____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__7____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__7____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[7].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__7____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__7____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__7____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__7____src_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[7].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__7____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__7____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__7____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__7____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[7].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__7____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__7____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__7____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__7____inc_src(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[7].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__7____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__6____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__6____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__6____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[6].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__6____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__6____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__6____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__6____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[6].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__6____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__6____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__6____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__6____src_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[6].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__6____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__6____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__6____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__6____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[6].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__6____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__6____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__6____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__6____inc_src(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[6].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__6____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__5____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__5____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__5____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[5].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__5____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__5____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__5____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__5____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[5].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__5____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__5____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__5____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__5____src_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[5].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__5____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__5____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__5____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__5____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[5].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__5____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__5____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__5____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__5____inc_src(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[5].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__5____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__4____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__4____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__4____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[4].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__4____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__4____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__4____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__4____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[4].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__4____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__4____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__4____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__4____src_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[4].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__4____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__4____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__4____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__4____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[4].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__4____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__4____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__4____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__4____inc_src(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[4].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__4____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__3____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__3____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__3____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[3].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__3____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__3____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__3____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__3____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[3].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__3____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__3____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__3____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__3____src_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[3].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__3____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__3____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__3____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__3____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[3].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__3____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__3____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__3____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__3____inc_src(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[3].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__3____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__2____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__2____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__2____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[2].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__2____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__2____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__2____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__2____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[2].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__2____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__2____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__2____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__2____src_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[2].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__2____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__2____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__2____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__2____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[2].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__2____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__2____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__2____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__2____inc_src(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[2].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__2____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__1____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__1____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__1____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[1].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__1____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__1____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__1____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__1____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[1].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__1____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__1____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__1____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__1____src_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[1].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__1____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__1____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__1____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__1____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[1].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__1____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__1____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__1____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__1____inc_src(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[1].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__1____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__0____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__0____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__0____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[0].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__0____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__0____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__0____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__0____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[0].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__0____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__0____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__0____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__0____src_sel(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[0].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__0____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__0____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__0____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__0____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[0].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__0____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t3__ll_desc__0____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__ll_desc__0____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t3__ll_desc__0____inc_src(longint unsigned meta_val);
        m_xfer_4par.t3.ll_desc[0].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__ll_desc__0____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t3__chk_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__chk_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t3__chk_sz(longint unsigned meta_val);
        m_xfer_4par.t3.chk_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__chk_sz::()>
//<unsigned_meta_action::_xfer_4par__t3__tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t3__tot_sz(longint unsigned meta_val);
        m_xfer_4par.t3.tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t3__dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__dst_sel(longint unsigned meta_val);
        m_xfer_4par.t3.dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__src_sel(longint unsigned meta_val);
        m_xfer_4par.t3.src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__src_sel::()>
//<unsigned_meta_action::_xfer_4par__t3__inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t3__inc_dst(longint unsigned meta_val);
        m_xfer_4par.t3.inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t3__inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t3__inc_src(longint unsigned meta_val);
        m_xfer_4par.t3.inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__inc_src::()>
//<unsigned_meta_action::_xfer_4par__t3__mode::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__mode
    //**************************************************************** 
   virtual task action_xfer_4par__t3__mode(longint unsigned meta_val);
        m_xfer_4par.t3.mode = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__mode::()>
//<unsigned_meta_action::_xfer_4par__t3__channel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t3__channel
    //**************************************************************** 
   virtual task action_xfer_4par__t3__channel(longint unsigned meta_val);
        m_xfer_4par.t3.channel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t3__channel::()>
//<unsigned_meta_action::_xfer_4par__t2__transfer_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__transfer_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t2__transfer_sz(longint unsigned meta_val);
        m_xfer_4par.t2.transfer_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__transfer_sz::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__15__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc_tot_sz__15__
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc_tot_sz__15__(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc_tot_sz[15] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__15__::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__14__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc_tot_sz__14__
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc_tot_sz__14__(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc_tot_sz[14] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__14__::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__13__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc_tot_sz__13__
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc_tot_sz__13__(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc_tot_sz[13] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__13__::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__12__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc_tot_sz__12__
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc_tot_sz__12__(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc_tot_sz[12] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__12__::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__11__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc_tot_sz__11__
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc_tot_sz__11__(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc_tot_sz[11] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__11__::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__10__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc_tot_sz__10__
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc_tot_sz__10__(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc_tot_sz[10] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__10__::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__9__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc_tot_sz__9__
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc_tot_sz__9__(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc_tot_sz[9] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__9__::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__8__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc_tot_sz__8__
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc_tot_sz__8__(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc_tot_sz[8] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__8__::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__7__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc_tot_sz__7__
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc_tot_sz__7__(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc_tot_sz[7] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__7__::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__6__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc_tot_sz__6__
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc_tot_sz__6__(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc_tot_sz[6] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__6__::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__5__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc_tot_sz__5__
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc_tot_sz__5__(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc_tot_sz[5] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__5__::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__4__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc_tot_sz__4__
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc_tot_sz__4__(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc_tot_sz[4] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__4__::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__3__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc_tot_sz__3__
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc_tot_sz__3__(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc_tot_sz[3] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__3__::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__2__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc_tot_sz__2__
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc_tot_sz__2__(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc_tot_sz[2] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__2__::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__1__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc_tot_sz__1__
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc_tot_sz__1__(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc_tot_sz[1] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__1__::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__0__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc_tot_sz__0__
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc_tot_sz__0__(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc_tot_sz[0] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc_tot_sz__0__::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc_sz(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc_sz::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__15____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__15____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__15____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[15].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__15____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__15____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__15____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__15____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[15].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__15____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__15____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__15____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__15____src_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[15].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__15____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__15____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__15____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__15____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[15].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__15____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__15____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__15____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__15____inc_src(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[15].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__15____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__14____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__14____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__14____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[14].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__14____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__14____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__14____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__14____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[14].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__14____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__14____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__14____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__14____src_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[14].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__14____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__14____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__14____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__14____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[14].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__14____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__14____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__14____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__14____inc_src(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[14].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__14____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__13____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__13____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__13____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[13].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__13____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__13____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__13____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__13____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[13].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__13____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__13____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__13____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__13____src_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[13].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__13____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__13____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__13____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__13____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[13].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__13____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__13____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__13____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__13____inc_src(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[13].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__13____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__12____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__12____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__12____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[12].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__12____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__12____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__12____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__12____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[12].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__12____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__12____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__12____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__12____src_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[12].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__12____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__12____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__12____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__12____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[12].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__12____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__12____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__12____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__12____inc_src(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[12].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__12____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__11____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__11____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__11____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[11].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__11____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__11____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__11____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__11____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[11].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__11____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__11____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__11____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__11____src_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[11].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__11____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__11____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__11____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__11____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[11].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__11____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__11____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__11____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__11____inc_src(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[11].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__11____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__10____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__10____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__10____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[10].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__10____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__10____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__10____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__10____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[10].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__10____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__10____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__10____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__10____src_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[10].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__10____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__10____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__10____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__10____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[10].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__10____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__10____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__10____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__10____inc_src(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[10].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__10____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__9____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__9____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__9____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[9].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__9____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__9____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__9____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__9____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[9].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__9____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__9____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__9____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__9____src_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[9].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__9____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__9____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__9____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__9____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[9].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__9____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__9____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__9____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__9____inc_src(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[9].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__9____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__8____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__8____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__8____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[8].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__8____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__8____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__8____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__8____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[8].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__8____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__8____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__8____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__8____src_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[8].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__8____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__8____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__8____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__8____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[8].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__8____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__8____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__8____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__8____inc_src(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[8].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__8____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__7____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__7____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__7____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[7].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__7____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__7____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__7____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__7____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[7].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__7____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__7____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__7____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__7____src_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[7].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__7____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__7____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__7____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__7____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[7].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__7____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__7____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__7____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__7____inc_src(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[7].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__7____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__6____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__6____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__6____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[6].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__6____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__6____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__6____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__6____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[6].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__6____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__6____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__6____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__6____src_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[6].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__6____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__6____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__6____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__6____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[6].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__6____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__6____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__6____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__6____inc_src(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[6].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__6____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__5____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__5____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__5____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[5].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__5____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__5____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__5____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__5____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[5].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__5____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__5____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__5____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__5____src_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[5].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__5____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__5____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__5____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__5____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[5].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__5____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__5____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__5____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__5____inc_src(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[5].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__5____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__4____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__4____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__4____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[4].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__4____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__4____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__4____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__4____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[4].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__4____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__4____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__4____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__4____src_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[4].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__4____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__4____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__4____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__4____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[4].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__4____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__4____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__4____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__4____inc_src(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[4].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__4____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__3____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__3____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__3____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[3].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__3____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__3____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__3____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__3____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[3].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__3____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__3____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__3____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__3____src_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[3].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__3____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__3____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__3____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__3____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[3].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__3____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__3____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__3____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__3____inc_src(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[3].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__3____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__2____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__2____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__2____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[2].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__2____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__2____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__2____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__2____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[2].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__2____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__2____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__2____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__2____src_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[2].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__2____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__2____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__2____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__2____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[2].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__2____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__2____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__2____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__2____inc_src(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[2].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__2____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__1____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__1____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__1____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[1].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__1____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__1____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__1____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__1____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[1].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__1____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__1____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__1____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__1____src_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[1].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__1____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__1____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__1____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__1____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[1].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__1____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__1____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__1____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__1____inc_src(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[1].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__1____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__0____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__0____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__0____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[0].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__0____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__0____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__0____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__0____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[0].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__0____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__0____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__0____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__0____src_sel(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[0].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__0____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__0____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__0____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__0____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[0].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__0____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t2__ll_desc__0____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__ll_desc__0____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t2__ll_desc__0____inc_src(longint unsigned meta_val);
        m_xfer_4par.t2.ll_desc[0].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__ll_desc__0____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t2__chk_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__chk_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t2__chk_sz(longint unsigned meta_val);
        m_xfer_4par.t2.chk_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__chk_sz::()>
//<unsigned_meta_action::_xfer_4par__t2__tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t2__tot_sz(longint unsigned meta_val);
        m_xfer_4par.t2.tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t2__dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__dst_sel(longint unsigned meta_val);
        m_xfer_4par.t2.dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__src_sel(longint unsigned meta_val);
        m_xfer_4par.t2.src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__src_sel::()>
//<unsigned_meta_action::_xfer_4par__t2__inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t2__inc_dst(longint unsigned meta_val);
        m_xfer_4par.t2.inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t2__inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t2__inc_src(longint unsigned meta_val);
        m_xfer_4par.t2.inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__inc_src::()>
//<unsigned_meta_action::_xfer_4par__t2__mode::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__mode
    //**************************************************************** 
   virtual task action_xfer_4par__t2__mode(longint unsigned meta_val);
        m_xfer_4par.t2.mode = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__mode::()>
//<unsigned_meta_action::_xfer_4par__t2__channel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t2__channel
    //**************************************************************** 
   virtual task action_xfer_4par__t2__channel(longint unsigned meta_val);
        m_xfer_4par.t2.channel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t2__channel::()>
//<unsigned_meta_action::_xfer_4par__t1__transfer_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__transfer_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t1__transfer_sz(longint unsigned meta_val);
        m_xfer_4par.t1.transfer_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__transfer_sz::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__15__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc_tot_sz__15__
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc_tot_sz__15__(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc_tot_sz[15] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__15__::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__14__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc_tot_sz__14__
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc_tot_sz__14__(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc_tot_sz[14] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__14__::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__13__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc_tot_sz__13__
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc_tot_sz__13__(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc_tot_sz[13] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__13__::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__12__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc_tot_sz__12__
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc_tot_sz__12__(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc_tot_sz[12] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__12__::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__11__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc_tot_sz__11__
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc_tot_sz__11__(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc_tot_sz[11] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__11__::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__10__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc_tot_sz__10__
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc_tot_sz__10__(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc_tot_sz[10] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__10__::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__9__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc_tot_sz__9__
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc_tot_sz__9__(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc_tot_sz[9] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__9__::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__8__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc_tot_sz__8__
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc_tot_sz__8__(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc_tot_sz[8] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__8__::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__7__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc_tot_sz__7__
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc_tot_sz__7__(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc_tot_sz[7] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__7__::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__6__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc_tot_sz__6__
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc_tot_sz__6__(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc_tot_sz[6] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__6__::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__5__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc_tot_sz__5__
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc_tot_sz__5__(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc_tot_sz[5] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__5__::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__4__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc_tot_sz__4__
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc_tot_sz__4__(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc_tot_sz[4] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__4__::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__3__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc_tot_sz__3__
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc_tot_sz__3__(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc_tot_sz[3] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__3__::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__2__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc_tot_sz__2__
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc_tot_sz__2__(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc_tot_sz[2] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__2__::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__1__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc_tot_sz__1__
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc_tot_sz__1__(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc_tot_sz[1] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__1__::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__0__::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc_tot_sz__0__
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc_tot_sz__0__(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc_tot_sz[0] = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc_tot_sz__0__::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc_sz(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc_sz::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__15____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__15____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__15____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[15].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__15____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__15____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__15____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__15____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[15].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__15____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__15____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__15____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__15____src_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[15].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__15____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__15____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__15____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__15____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[15].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__15____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__15____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__15____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__15____inc_src(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[15].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__15____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__14____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__14____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__14____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[14].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__14____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__14____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__14____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__14____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[14].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__14____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__14____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__14____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__14____src_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[14].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__14____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__14____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__14____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__14____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[14].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__14____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__14____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__14____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__14____inc_src(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[14].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__14____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__13____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__13____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__13____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[13].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__13____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__13____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__13____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__13____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[13].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__13____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__13____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__13____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__13____src_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[13].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__13____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__13____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__13____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__13____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[13].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__13____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__13____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__13____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__13____inc_src(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[13].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__13____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__12____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__12____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__12____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[12].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__12____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__12____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__12____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__12____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[12].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__12____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__12____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__12____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__12____src_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[12].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__12____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__12____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__12____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__12____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[12].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__12____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__12____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__12____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__12____inc_src(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[12].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__12____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__11____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__11____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__11____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[11].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__11____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__11____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__11____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__11____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[11].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__11____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__11____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__11____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__11____src_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[11].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__11____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__11____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__11____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__11____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[11].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__11____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__11____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__11____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__11____inc_src(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[11].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__11____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__10____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__10____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__10____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[10].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__10____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__10____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__10____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__10____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[10].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__10____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__10____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__10____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__10____src_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[10].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__10____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__10____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__10____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__10____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[10].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__10____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__10____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__10____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__10____inc_src(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[10].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__10____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__9____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__9____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__9____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[9].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__9____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__9____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__9____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__9____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[9].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__9____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__9____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__9____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__9____src_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[9].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__9____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__9____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__9____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__9____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[9].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__9____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__9____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__9____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__9____inc_src(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[9].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__9____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__8____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__8____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__8____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[8].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__8____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__8____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__8____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__8____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[8].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__8____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__8____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__8____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__8____src_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[8].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__8____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__8____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__8____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__8____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[8].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__8____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__8____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__8____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__8____inc_src(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[8].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__8____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__7____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__7____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__7____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[7].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__7____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__7____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__7____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__7____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[7].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__7____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__7____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__7____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__7____src_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[7].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__7____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__7____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__7____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__7____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[7].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__7____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__7____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__7____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__7____inc_src(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[7].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__7____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__6____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__6____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__6____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[6].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__6____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__6____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__6____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__6____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[6].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__6____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__6____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__6____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__6____src_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[6].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__6____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__6____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__6____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__6____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[6].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__6____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__6____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__6____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__6____inc_src(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[6].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__6____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__5____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__5____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__5____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[5].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__5____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__5____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__5____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__5____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[5].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__5____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__5____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__5____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__5____src_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[5].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__5____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__5____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__5____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__5____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[5].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__5____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__5____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__5____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__5____inc_src(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[5].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__5____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__4____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__4____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__4____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[4].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__4____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__4____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__4____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__4____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[4].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__4____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__4____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__4____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__4____src_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[4].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__4____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__4____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__4____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__4____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[4].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__4____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__4____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__4____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__4____inc_src(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[4].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__4____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__3____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__3____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__3____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[3].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__3____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__3____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__3____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__3____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[3].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__3____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__3____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__3____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__3____src_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[3].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__3____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__3____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__3____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__3____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[3].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__3____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__3____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__3____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__3____inc_src(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[3].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__3____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__2____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__2____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__2____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[2].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__2____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__2____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__2____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__2____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[2].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__2____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__2____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__2____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__2____src_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[2].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__2____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__2____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__2____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__2____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[2].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__2____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__2____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__2____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__2____inc_src(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[2].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__2____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__1____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__1____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__1____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[1].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__1____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__1____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__1____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__1____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[1].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__1____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__1____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__1____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__1____src_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[1].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__1____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__1____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__1____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__1____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[1].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__1____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__1____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__1____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__1____inc_src(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[1].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__1____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__0____tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__0____tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__0____tot_sz(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[0].tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__0____tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__0____dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__0____dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__0____dst_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[0].dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__0____dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__0____src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__0____src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__0____src_sel(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[0].src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__0____src_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__0____inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__0____inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__0____inc_dst(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[0].inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__0____inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t1__ll_desc__0____inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__ll_desc__0____inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t1__ll_desc__0____inc_src(longint unsigned meta_val);
        m_xfer_4par.t1.ll_desc[0].inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__ll_desc__0____inc_src::()>
//<unsigned_meta_action::_xfer_4par__t1__chk_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__chk_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t1__chk_sz(longint unsigned meta_val);
        m_xfer_4par.t1.chk_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__chk_sz::()>
//<unsigned_meta_action::_xfer_4par__t1__tot_sz::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__tot_sz
    //**************************************************************** 
   virtual task action_xfer_4par__t1__tot_sz(longint unsigned meta_val);
        m_xfer_4par.t1.tot_sz = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__tot_sz::()>
//<unsigned_meta_action::_xfer_4par__t1__dst_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__dst_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__dst_sel(longint unsigned meta_val);
        m_xfer_4par.t1.dst_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__dst_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__src_sel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__src_sel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__src_sel(longint unsigned meta_val);
        m_xfer_4par.t1.src_sel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__src_sel::()>
//<unsigned_meta_action::_xfer_4par__t1__inc_dst::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__inc_dst
    //**************************************************************** 
   virtual task action_xfer_4par__t1__inc_dst(longint unsigned meta_val);
        m_xfer_4par.t1.inc_dst = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__inc_dst::()>
//<unsigned_meta_action::_xfer_4par__t1__inc_src::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__inc_src
    //**************************************************************** 
   virtual task action_xfer_4par__t1__inc_src(longint unsigned meta_val);
        m_xfer_4par.t1.inc_src = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__inc_src::()>
//<unsigned_meta_action::_xfer_4par__t1__mode::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__mode
    //**************************************************************** 
   virtual task action_xfer_4par__t1__mode(longint unsigned meta_val);
        m_xfer_4par.t1.mode = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__mode::()>
//<unsigned_meta_action::_xfer_4par__t1__channel::()>
    //***************************************************************
    //* Action task action_xfer_4par__t1__channel
    //**************************************************************** 
   virtual task action_xfer_4par__t1__channel(longint unsigned meta_val);
        m_xfer_4par.t1.channel = meta_val;
    endtask
//</unsigned_meta_action::_xfer_4par__t1__channel::()>
//<action::_wait_done::()>
    //***************************************************************
    //* Action task action_wait_done
    //**************************************************************** 
   virtual task action_wait_done();
    endtask
//</action::_wait_done::()>
//</trashcan>
`endif


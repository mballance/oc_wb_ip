
`include "uvm_macros.svh"

package wb_uart_env_pkg;
	import uvm_pkg::*;
	import wb_master_agent_pkg::*;

	`include "wb_uart_env.svh"
	
endpackage

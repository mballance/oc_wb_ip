/****************************************************************************
 * wb_mem_mgr.svh
 ****************************************************************************/

/**
 * Class: wb_mem_mgr
 * 
 * TODO: Add class documentation
 */
class wb_mem_mgr;

	function new();

	endfunction


endclass



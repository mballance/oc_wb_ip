
`include "uvm_macros.svh"

package wb_simple_pic_env_pkg;
	import uvm_pkg::*;

	`include "wb_simple_pic_env.svh"
	
endpackage

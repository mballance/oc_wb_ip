

`include "uvm_macros.svh"
package wb_periph_subsys_tests_pkg;
	import uvm_pkg::*;
	import wb_periph_subsys_env_pkg::*;
	
	`include "wb_periph_subsys_test_base.svh"
	
endpackage

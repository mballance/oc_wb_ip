
`include "uvm_macros.svh"

package wb_uart16550_env_pkg;
	import uvm_pkg::*;
	import wb_master_agent_pkg::*;
	import sv_bfms_api_pkg::*;

	`include "wb_uart16550_env.svh"
	
endpackage

/****************************************************************************
 * wb_periph_subsys_vseq.svh
 ****************************************************************************/

/**
 * Class: wb_periph_subsys_vseq
 * 
 * TODO: Add class documentation
 */
class wb_periph_subsys_vseq extends uvm_sequence;

	function new();

	endfunction


endclass



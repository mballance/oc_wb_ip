
`include "uvm_macros.svh"

package wb_dma_env_pkg;
	import uvm_pkg::*;
	import wb_dma_regs_pkg::*;

	`include "wb_dma_env.svh"
	
endpackage

/****************************************************************************
 * wb_dma_dev_pkg.sv
 ****************************************************************************/
`include "uvm_macros.svh"
`include "uvmdev_macros.svh"

/**
 * Package: wb_dma_dev_pkg
 * 
 * TODO: Add package documentation
 */
package wb_dma_dev_pkg;
	import uvm_pkg::*;
	import uvmdev_pkg::*;
	import wb_dma_regs_pkg::*;

	`include "wb_dma_dev.svh"
	
endpackage





`include "uvm_macros.svh"
package wb_simple_pic_tests_pkg;
	import uvm_pkg::*;
	import wb_simple_pic_env_pkg::*;
	
	`include "wb_simple_pic_test_base.svh"
	
endpackage


`line 1 "wb_dma_infact_4par_seq.svh" 0






   
`line 7 "wb_dma_infact_4par_seq.svh" 0

  
`line 8 "wb_dma_infact_4par_seq.svh" 0






  
`line 1 "wb_dma_infact_4par_seq_scheduler.svh" 0

`line 1 "wb_dma_infact_4par_seq_scheduler.svh" 0

        
           


  
`line 6 "wb_dma_infact_4par_seq_scheduler.svh" 0

  
`line 7 "wb_dma_infact_4par_seq_scheduler.svh" 0


import inFactSv::*;

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_infact_checkcov #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_actionTask(te, "infact_checkcov");
  endfunction
  task actionTask();
    _parent.action_infact_checkcov();
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_infact_checkcov

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_wait_done #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_actionTask(te, "wait_done");
  endfunction
  task actionTask();
    _parent.action_wait_done();
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_wait_done

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_init_xfer__t4__end #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_actionTask(te, "init_xfer(t4).end");
  endfunction
  task actionTask();
    _parent.action_init_xfer__t4__end();
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_init_xfer__t4__end

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_init_xfer__t4__begin #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_actionTask(te, "init_xfer(t4).begin");
  endfunction
  task actionTask();
    _parent.action_init_xfer__t4__begin();
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_init_xfer__t4__begin

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_init_xfer__t3__end #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_actionTask(te, "init_xfer(t3).end");
  endfunction
  task actionTask();
    _parent.action_init_xfer__t3__end();
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_init_xfer__t3__end

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_init_xfer__t3__begin #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_actionTask(te, "init_xfer(t3).begin");
  endfunction
  task actionTask();
    _parent.action_init_xfer__t3__begin();
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_init_xfer__t3__begin

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_init_xfer__t2__end #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_actionTask(te, "init_xfer(t2).end");
  endfunction
  task actionTask();
    _parent.action_init_xfer__t2__end();
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_init_xfer__t2__end

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_init_xfer__t2__begin #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_actionTask(te, "init_xfer(t2).begin");
  endfunction
  task actionTask();
    _parent.action_init_xfer__t2__begin();
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_init_xfer__t2__begin

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_init_xfer__t1__end #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_actionTask(te, "init_xfer(t1).end");
  endfunction
  task actionTask();
    _parent.action_init_xfer__t1__end();
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_init_xfer__t1__end

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_init_xfer__t1__begin #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_actionTask(te, "init_xfer(t1).begin");
  endfunction
  task actionTask();
    _parent.action_init_xfer__t1__begin();
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_init_xfer__t1__begin

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_init #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_actionTask(te, "init");
  endfunction
  task actionTask();
    _parent.action_init();
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_init

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__sum #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_signedMetaActionTask(te, "t4.ll_desc_tot_sz.sum");
  endfunction
  task signedMetaActionTask(input longint signed value);
    _parent.action_t4__ll_desc_tot_sz__sum(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__sum

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__sum #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_signedMetaActionTask(te, "t3.ll_desc_tot_sz.sum");
  endfunction
  task signedMetaActionTask(input longint signed value);
    _parent.action_t3__ll_desc_tot_sz__sum(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__sum

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__sum #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_signedMetaActionTask(te, "t2.ll_desc_tot_sz.sum");
  endfunction
  task signedMetaActionTask(input longint signed value);
    _parent.action_t2__ll_desc_tot_sz__sum(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__sum

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__sum #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_signedMetaActionTask(te, "t1.ll_desc_tot_sz.sum");
  endfunction
  task signedMetaActionTask(input longint signed value);
    _parent.action_t1__ll_desc_tot_sz__sum(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__sum

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__transfer_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.transfer_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__transfer_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__transfer_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__15__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc_tot_sz[15]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc_tot_sz__15__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__15__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__14__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc_tot_sz[14]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc_tot_sz__14__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__14__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__13__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc_tot_sz[13]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc_tot_sz__13__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__13__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__12__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc_tot_sz[12]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc_tot_sz__12__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__12__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__11__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc_tot_sz[11]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc_tot_sz__11__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__11__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__10__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc_tot_sz[10]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc_tot_sz__10__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__10__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__9__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc_tot_sz[9]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc_tot_sz__9__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__9__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__8__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc_tot_sz[8]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc_tot_sz__8__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__8__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__7__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc_tot_sz[7]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc_tot_sz__7__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__7__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__6__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc_tot_sz[6]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc_tot_sz__6__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__6__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__5__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc_tot_sz[5]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc_tot_sz__5__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__5__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__4__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc_tot_sz[4]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc_tot_sz__4__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__4__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__3__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc_tot_sz[3]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc_tot_sz__3__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__3__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__2__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc_tot_sz[2]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc_tot_sz__2__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__2__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__1__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc_tot_sz[1]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc_tot_sz__1__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__1__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__0__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc_tot_sz[0]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc_tot_sz__0__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_tot_sz__0__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__15____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[15].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__15____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__15____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__15____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[15].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__15____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__15____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__15____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[15].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__15____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__15____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__15____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[15].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__15____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__15____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__15____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[15].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__15____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__15____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__14____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[14].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__14____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__14____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__14____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[14].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__14____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__14____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__14____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[14].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__14____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__14____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__14____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[14].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__14____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__14____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__14____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[14].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__14____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__14____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__13____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[13].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__13____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__13____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__13____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[13].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__13____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__13____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__13____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[13].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__13____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__13____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__13____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[13].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__13____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__13____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__13____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[13].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__13____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__13____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__12____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[12].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__12____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__12____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__12____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[12].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__12____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__12____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__12____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[12].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__12____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__12____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__12____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[12].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__12____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__12____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__12____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[12].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__12____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__12____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__11____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[11].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__11____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__11____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__11____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[11].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__11____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__11____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__11____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[11].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__11____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__11____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__11____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[11].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__11____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__11____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__11____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[11].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__11____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__11____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__10____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[10].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__10____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__10____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__10____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[10].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__10____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__10____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__10____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[10].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__10____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__10____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__10____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[10].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__10____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__10____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__10____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[10].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__10____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__10____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__9____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[9].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__9____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__9____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__9____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[9].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__9____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__9____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__9____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[9].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__9____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__9____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__9____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[9].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__9____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__9____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__9____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[9].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__9____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__9____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__8____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[8].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__8____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__8____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__8____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[8].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__8____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__8____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__8____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[8].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__8____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__8____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__8____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[8].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__8____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__8____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__8____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[8].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__8____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__8____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__7____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[7].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__7____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__7____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__7____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[7].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__7____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__7____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__7____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[7].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__7____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__7____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__7____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[7].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__7____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__7____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__7____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[7].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__7____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__7____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__6____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[6].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__6____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__6____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__6____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[6].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__6____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__6____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__6____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[6].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__6____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__6____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__6____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[6].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__6____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__6____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__6____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[6].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__6____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__6____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__5____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[5].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__5____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__5____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__5____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[5].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__5____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__5____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__5____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[5].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__5____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__5____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__5____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[5].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__5____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__5____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__5____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[5].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__5____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__5____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__4____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[4].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__4____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__4____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__4____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[4].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__4____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__4____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__4____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[4].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__4____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__4____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__4____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[4].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__4____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__4____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__4____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[4].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__4____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__4____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__3____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[3].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__3____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__3____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__3____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[3].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__3____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__3____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__3____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[3].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__3____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__3____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__3____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[3].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__3____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__3____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__3____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[3].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__3____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__3____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__2____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[2].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__2____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__2____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__2____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[2].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__2____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__2____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__2____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[2].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__2____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__2____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__2____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[2].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__2____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__2____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__2____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[2].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__2____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__2____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__1____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[1].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__1____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__1____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__1____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[1].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__1____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__1____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__1____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[1].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__1____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__1____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__1____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[1].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__1____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__1____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__1____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[1].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__1____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__1____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__0____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[0].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__0____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__0____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__0____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[0].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__0____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__0____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__0____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[0].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__0____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__0____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__0____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[0].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__0____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__0____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__0____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.ll_desc[0].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__ll_desc__0____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__ll_desc__0____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__chk_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.chk_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__chk_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__chk_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__mode #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.mode");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__mode(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__mode

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__channel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t4.channel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t4__channel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t4__channel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__transfer_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.transfer_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__transfer_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__transfer_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__15__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc_tot_sz[15]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc_tot_sz__15__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__15__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__14__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc_tot_sz[14]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc_tot_sz__14__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__14__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__13__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc_tot_sz[13]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc_tot_sz__13__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__13__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__12__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc_tot_sz[12]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc_tot_sz__12__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__12__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__11__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc_tot_sz[11]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc_tot_sz__11__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__11__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__10__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc_tot_sz[10]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc_tot_sz__10__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__10__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__9__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc_tot_sz[9]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc_tot_sz__9__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__9__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__8__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc_tot_sz[8]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc_tot_sz__8__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__8__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__7__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc_tot_sz[7]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc_tot_sz__7__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__7__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__6__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc_tot_sz[6]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc_tot_sz__6__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__6__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__5__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc_tot_sz[5]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc_tot_sz__5__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__5__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__4__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc_tot_sz[4]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc_tot_sz__4__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__4__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__3__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc_tot_sz[3]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc_tot_sz__3__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__3__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__2__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc_tot_sz[2]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc_tot_sz__2__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__2__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__1__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc_tot_sz[1]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc_tot_sz__1__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__1__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__0__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc_tot_sz[0]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc_tot_sz__0__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_tot_sz__0__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__15____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[15].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__15____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__15____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__15____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[15].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__15____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__15____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__15____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[15].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__15____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__15____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__15____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[15].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__15____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__15____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__15____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[15].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__15____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__15____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__14____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[14].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__14____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__14____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__14____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[14].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__14____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__14____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__14____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[14].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__14____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__14____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__14____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[14].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__14____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__14____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__14____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[14].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__14____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__14____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__13____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[13].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__13____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__13____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__13____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[13].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__13____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__13____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__13____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[13].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__13____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__13____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__13____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[13].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__13____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__13____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__13____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[13].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__13____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__13____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__12____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[12].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__12____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__12____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__12____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[12].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__12____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__12____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__12____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[12].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__12____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__12____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__12____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[12].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__12____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__12____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__12____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[12].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__12____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__12____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__11____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[11].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__11____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__11____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__11____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[11].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__11____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__11____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__11____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[11].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__11____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__11____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__11____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[11].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__11____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__11____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__11____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[11].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__11____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__11____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__10____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[10].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__10____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__10____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__10____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[10].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__10____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__10____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__10____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[10].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__10____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__10____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__10____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[10].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__10____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__10____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__10____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[10].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__10____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__10____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__9____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[9].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__9____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__9____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__9____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[9].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__9____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__9____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__9____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[9].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__9____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__9____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__9____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[9].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__9____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__9____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__9____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[9].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__9____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__9____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__8____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[8].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__8____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__8____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__8____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[8].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__8____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__8____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__8____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[8].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__8____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__8____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__8____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[8].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__8____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__8____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__8____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[8].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__8____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__8____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__7____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[7].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__7____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__7____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__7____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[7].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__7____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__7____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__7____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[7].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__7____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__7____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__7____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[7].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__7____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__7____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__7____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[7].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__7____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__7____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__6____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[6].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__6____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__6____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__6____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[6].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__6____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__6____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__6____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[6].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__6____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__6____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__6____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[6].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__6____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__6____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__6____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[6].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__6____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__6____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__5____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[5].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__5____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__5____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__5____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[5].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__5____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__5____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__5____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[5].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__5____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__5____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__5____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[5].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__5____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__5____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__5____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[5].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__5____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__5____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__4____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[4].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__4____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__4____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__4____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[4].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__4____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__4____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__4____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[4].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__4____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__4____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__4____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[4].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__4____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__4____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__4____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[4].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__4____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__4____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__3____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[3].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__3____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__3____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__3____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[3].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__3____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__3____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__3____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[3].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__3____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__3____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__3____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[3].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__3____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__3____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__3____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[3].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__3____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__3____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__2____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[2].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__2____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__2____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__2____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[2].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__2____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__2____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__2____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[2].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__2____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__2____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__2____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[2].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__2____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__2____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__2____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[2].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__2____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__2____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__1____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[1].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__1____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__1____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__1____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[1].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__1____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__1____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__1____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[1].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__1____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__1____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__1____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[1].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__1____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__1____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__1____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[1].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__1____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__1____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__0____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[0].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__0____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__0____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__0____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[0].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__0____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__0____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__0____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[0].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__0____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__0____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__0____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[0].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__0____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__0____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__0____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.ll_desc[0].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__ll_desc__0____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__ll_desc__0____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__chk_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.chk_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__chk_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__chk_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__mode #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.mode");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__mode(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__mode

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__channel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t3.channel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t3__channel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t3__channel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__transfer_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.transfer_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__transfer_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__transfer_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__15__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc_tot_sz[15]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc_tot_sz__15__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__15__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__14__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc_tot_sz[14]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc_tot_sz__14__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__14__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__13__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc_tot_sz[13]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc_tot_sz__13__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__13__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__12__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc_tot_sz[12]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc_tot_sz__12__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__12__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__11__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc_tot_sz[11]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc_tot_sz__11__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__11__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__10__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc_tot_sz[10]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc_tot_sz__10__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__10__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__9__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc_tot_sz[9]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc_tot_sz__9__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__9__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__8__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc_tot_sz[8]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc_tot_sz__8__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__8__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__7__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc_tot_sz[7]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc_tot_sz__7__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__7__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__6__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc_tot_sz[6]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc_tot_sz__6__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__6__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__5__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc_tot_sz[5]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc_tot_sz__5__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__5__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__4__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc_tot_sz[4]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc_tot_sz__4__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__4__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__3__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc_tot_sz[3]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc_tot_sz__3__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__3__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__2__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc_tot_sz[2]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc_tot_sz__2__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__2__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__1__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc_tot_sz[1]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc_tot_sz__1__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__1__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__0__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc_tot_sz[0]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc_tot_sz__0__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_tot_sz__0__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__15____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[15].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__15____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__15____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__15____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[15].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__15____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__15____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__15____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[15].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__15____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__15____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__15____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[15].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__15____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__15____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__15____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[15].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__15____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__15____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__14____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[14].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__14____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__14____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__14____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[14].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__14____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__14____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__14____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[14].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__14____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__14____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__14____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[14].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__14____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__14____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__14____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[14].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__14____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__14____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__13____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[13].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__13____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__13____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__13____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[13].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__13____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__13____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__13____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[13].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__13____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__13____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__13____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[13].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__13____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__13____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__13____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[13].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__13____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__13____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__12____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[12].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__12____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__12____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__12____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[12].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__12____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__12____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__12____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[12].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__12____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__12____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__12____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[12].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__12____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__12____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__12____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[12].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__12____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__12____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__11____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[11].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__11____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__11____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__11____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[11].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__11____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__11____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__11____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[11].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__11____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__11____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__11____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[11].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__11____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__11____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__11____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[11].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__11____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__11____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__10____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[10].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__10____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__10____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__10____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[10].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__10____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__10____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__10____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[10].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__10____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__10____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__10____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[10].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__10____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__10____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__10____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[10].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__10____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__10____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__9____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[9].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__9____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__9____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__9____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[9].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__9____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__9____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__9____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[9].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__9____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__9____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__9____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[9].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__9____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__9____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__9____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[9].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__9____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__9____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__8____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[8].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__8____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__8____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__8____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[8].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__8____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__8____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__8____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[8].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__8____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__8____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__8____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[8].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__8____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__8____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__8____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[8].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__8____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__8____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__7____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[7].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__7____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__7____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__7____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[7].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__7____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__7____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__7____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[7].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__7____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__7____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__7____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[7].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__7____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__7____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__7____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[7].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__7____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__7____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__6____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[6].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__6____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__6____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__6____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[6].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__6____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__6____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__6____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[6].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__6____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__6____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__6____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[6].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__6____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__6____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__6____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[6].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__6____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__6____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__5____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[5].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__5____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__5____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__5____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[5].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__5____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__5____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__5____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[5].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__5____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__5____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__5____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[5].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__5____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__5____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__5____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[5].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__5____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__5____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__4____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[4].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__4____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__4____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__4____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[4].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__4____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__4____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__4____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[4].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__4____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__4____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__4____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[4].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__4____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__4____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__4____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[4].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__4____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__4____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__3____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[3].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__3____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__3____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__3____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[3].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__3____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__3____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__3____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[3].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__3____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__3____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__3____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[3].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__3____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__3____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__3____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[3].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__3____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__3____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__2____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[2].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__2____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__2____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__2____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[2].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__2____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__2____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__2____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[2].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__2____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__2____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__2____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[2].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__2____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__2____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__2____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[2].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__2____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__2____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__1____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[1].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__1____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__1____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__1____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[1].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__1____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__1____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__1____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[1].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__1____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__1____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__1____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[1].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__1____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__1____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__1____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[1].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__1____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__1____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__0____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[0].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__0____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__0____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__0____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[0].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__0____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__0____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__0____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[0].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__0____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__0____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__0____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[0].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__0____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__0____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__0____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.ll_desc[0].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__ll_desc__0____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__ll_desc__0____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__chk_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.chk_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__chk_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__chk_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__mode #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.mode");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__mode(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__mode

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__channel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t2.channel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t2__channel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t2__channel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__transfer_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.transfer_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__transfer_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__transfer_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__15__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc_tot_sz[15]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc_tot_sz__15__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__15__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__14__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc_tot_sz[14]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc_tot_sz__14__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__14__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__13__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc_tot_sz[13]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc_tot_sz__13__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__13__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__12__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc_tot_sz[12]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc_tot_sz__12__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__12__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__11__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc_tot_sz[11]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc_tot_sz__11__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__11__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__10__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc_tot_sz[10]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc_tot_sz__10__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__10__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__9__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc_tot_sz[9]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc_tot_sz__9__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__9__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__8__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc_tot_sz[8]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc_tot_sz__8__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__8__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__7__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc_tot_sz[7]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc_tot_sz__7__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__7__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__6__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc_tot_sz[6]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc_tot_sz__6__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__6__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__5__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc_tot_sz[5]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc_tot_sz__5__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__5__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__4__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc_tot_sz[4]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc_tot_sz__4__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__4__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__3__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc_tot_sz[3]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc_tot_sz__3__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__3__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__2__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc_tot_sz[2]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc_tot_sz__2__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__2__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__1__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc_tot_sz[1]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc_tot_sz__1__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__1__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__0__ #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc_tot_sz[0]");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc_tot_sz__0__(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_tot_sz__0__

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__15____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[15].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__15____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__15____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__15____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[15].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__15____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__15____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__15____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[15].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__15____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__15____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__15____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[15].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__15____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__15____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__15____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[15].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__15____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__15____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__14____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[14].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__14____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__14____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__14____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[14].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__14____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__14____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__14____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[14].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__14____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__14____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__14____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[14].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__14____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__14____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__14____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[14].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__14____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__14____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__13____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[13].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__13____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__13____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__13____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[13].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__13____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__13____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__13____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[13].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__13____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__13____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__13____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[13].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__13____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__13____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__13____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[13].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__13____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__13____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__12____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[12].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__12____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__12____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__12____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[12].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__12____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__12____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__12____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[12].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__12____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__12____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__12____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[12].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__12____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__12____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__12____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[12].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__12____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__12____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__11____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[11].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__11____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__11____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__11____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[11].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__11____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__11____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__11____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[11].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__11____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__11____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__11____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[11].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__11____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__11____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__11____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[11].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__11____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__11____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__10____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[10].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__10____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__10____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__10____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[10].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__10____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__10____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__10____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[10].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__10____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__10____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__10____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[10].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__10____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__10____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__10____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[10].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__10____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__10____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__9____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[9].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__9____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__9____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__9____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[9].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__9____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__9____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__9____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[9].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__9____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__9____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__9____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[9].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__9____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__9____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__9____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[9].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__9____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__9____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__8____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[8].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__8____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__8____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__8____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[8].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__8____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__8____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__8____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[8].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__8____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__8____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__8____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[8].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__8____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__8____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__8____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[8].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__8____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__8____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__7____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[7].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__7____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__7____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__7____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[7].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__7____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__7____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__7____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[7].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__7____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__7____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__7____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[7].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__7____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__7____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__7____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[7].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__7____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__7____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__6____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[6].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__6____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__6____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__6____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[6].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__6____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__6____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__6____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[6].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__6____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__6____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__6____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[6].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__6____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__6____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__6____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[6].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__6____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__6____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__5____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[5].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__5____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__5____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__5____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[5].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__5____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__5____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__5____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[5].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__5____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__5____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__5____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[5].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__5____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__5____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__5____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[5].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__5____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__5____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__4____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[4].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__4____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__4____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__4____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[4].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__4____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__4____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__4____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[4].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__4____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__4____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__4____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[4].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__4____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__4____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__4____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[4].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__4____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__4____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__3____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[3].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__3____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__3____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__3____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[3].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__3____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__3____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__3____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[3].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__3____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__3____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__3____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[3].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__3____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__3____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__3____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[3].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__3____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__3____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__2____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[2].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__2____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__2____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__2____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[2].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__2____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__2____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__2____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[2].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__2____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__2____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__2____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[2].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__2____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__2____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__2____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[2].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__2____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__2____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__1____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[1].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__1____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__1____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__1____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[1].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__1____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__1____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__1____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[1].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__1____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__1____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__1____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[1].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__1____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__1____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__1____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[1].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__1____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__1____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__0____tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[0].tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__0____tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__0____tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__0____dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[0].dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__0____dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__0____dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__0____src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[0].src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__0____src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__0____src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__0____inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[0].inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__0____inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__0____inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__0____inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.ll_desc[0].inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__ll_desc__0____inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__ll_desc__0____inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__chk_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.chk_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__chk_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__chk_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__tot_sz #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.tot_sz");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__tot_sz(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__tot_sz

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__dst_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.dst_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__dst_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__dst_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__src_sel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.src_sel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__src_sel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__src_sel

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__inc_dst #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.inc_dst");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__inc_dst(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__inc_dst

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__inc_src #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.inc_src");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__inc_src(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__inc_src

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__mode #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.mode");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__mode(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__mode

class wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__channel #(type T=int) extends inFactSv::FunctorBase;
  T _parent;
  inFactSv::TestEngine thisTestEngine;
  function new(T parent, inFactSv::TestEngine te);
    _parent = parent;
    thisTestEngine = te;
    register_unsignedMetaActionTask(te, "t1.channel");
  endfunction
  task unsignedMetaActionTask(input longint unsigned value);
    _parent.action_t1__channel(value);
  endtask
endclass: wb_dma_infact_4par_seq_scheduler_wb_dma_infact_4par_seq_t1__channel

class wb_dma_infact_4par_seq_scheduler;
  inFactSv::TestEngine _wb_dma_infact_4par_seq_te;
  function new(string instanceName);
    _wb_dma_infact_4par_seq_te = new($psprintf("wb_dma_infact_4par_seq()"), instanceName, "wb_dma_infact_4par_seq_scheduler", 1, 0, $psprintf(""));
  endfunction
  task run_all();
    fork
      run_wb_dma_infact_4par_seq();
    join
  endtask: run_all
  task run_wb_dma_infact_4par_seq();
    _wb_dma_infact_4par_seq_te.run();
  endtask: run_wb_dma_infact_4par_seq
  task suspend_immediately_wb_dma_infact_4par_seq();
    disable run_wb_dma_infact_4par_seq;
  endtask: suspend_immediately_wb_dma_infact_4par_seq
  function inFactSv::TestEngine wb_dma_infact_4par_seq();
    return _wb_dma_infact_4par_seq_te;
  endfunction
endclass: wb_dma_infact_4par_seq_scheduler

 
`line 5739 "wb_dma_infact_4par_seq_scheduler.svh" 0
 

`line 5740 "wb_dma_infact_4par_seq.svh" 0



  
`line 1 "wb_dma_infact_4par_seq_items.svh" 0

`line 1 "wb_dma_infact_4par_seq_items.svh" 0

 

      

  
`line 6 "wb_dma_infact_4par_seq_items.svh" 0

  
`line 7 "wb_dma_infact_4par_seq_items.svh" 0


class wb_dma_infact_4par_seq_enums_c;
endclass


class wb_dma_infact_4par_seq_uvm_void_c;
endclass


class wb_dma_infact_4par_seq_uvm_object_c extends wb_dma_infact_4par_seq_uvm_void_c;
endclass


class wb_dma_infact_4par_seq_wb_dma_ll_descriptor_c extends wb_dma_infact_4par_seq_uvm_object_c;
    bit[63:0]		inc_src;
    bit[63:0]		inc_dst;
    bit[63:0]		src_sel;
    bit[63:0]		dst_sel;
    bit[63:0]		tot_sz;
endclass


class wb_dma_infact_4par_seq_wb_dma_descriptor_c;
    bit[63:0]		channel;
    bit[63:0]		mode;
    bit[63:0]		inc_src;
    bit[63:0]		inc_dst;
    bit[63:0]		src_sel;
    bit[63:0]		dst_sel;
    bit[63:0]		tot_sz;
    bit[63:0]		chk_sz;
    wb_dma_infact_4par_seq_wb_dma_ll_descriptor_c		ll_desc[16];
    bit[63:0]		ll_desc_sz;
    bit[63:0]		ll_desc_tot_sz[16];
    bit signed [63:0]		ll_desc_tot_sz__sum;
    bit[63:0]		transfer_sz;

    function new();
        for (int index__0 = 0; index__0 < 16; index__0++)
            ll_desc[index__0] = new();
    endfunction
endclass






 
`line 56 "wb_dma_infact_4par_seq_items.svh" 0
  


`line 58 "wb_dma_infact_4par_seq.svh" 0


  
`line 1 "wb_dma_infact_4par_seq_fields_cov.svh" 0

`line 1 "wb_dma_infact_4par_seq_fields_cov.svh" 0

 

        

       

  
`line 8 "wb_dma_infact_4par_seq_fields_cov.svh" 0

  
`line 9 "wb_dma_infact_4par_seq_fields_cov.svh" 0




class wb_dma_infact_4par_seq_fields_cov;

	
	
	
    PathCoverage              m_t1_channel_ac;
    PathCoverage              m_t2_channel_ac;
    PathCoverage              m_t3_channel_ac;
    PathCoverage              m_t4_channel_ac;


	
	PathCoverage						m_path_coverages[$];
	
	string								m_inst_name;

	

	
 

    

	function new(TestEngine eng, string inst_name="", bit instantiate_fc=1);
		string basename = inst_name;
		if (inst_name != "") begin
			inst_name = {inst_name, "."};
			m_inst_name = inst_name;
		end else begin
			m_inst_name = "";
		end
		
		if (instantiate_fc) begin

		end
        
        m_t1_channel_ac = new("t1.channel", {inst_name, "t1_channel_ac"}, eng);
        m_t1_channel_ac.addPathStopNode("t1.channel");
        m_t1_channel_ac.setGoalPathHitCount(1);
        m_t1_channel_ac.addBinScheme("wb_dma_infact_4par_seq_fields_cov_bin_scheme");
        m_t1_channel_ac.addPathConstraint("wb_dma_infact_4par_seq_fields_cov_bin_scheme$__unbinned_filter");
        m_t1_channel_ac.setSpecificationComplete();
        m_path_coverages.push_back(m_t1_channel_ac);


        
        m_t2_channel_ac = new("t2.channel", {inst_name, "t2_channel_ac"}, eng);
        m_t2_channel_ac.addPathStopNode("t2.channel");
        m_t2_channel_ac.setGoalPathHitCount(1);
        m_t2_channel_ac.addBinScheme("wb_dma_infact_4par_seq_fields_cov_bin_scheme");
        m_t2_channel_ac.addPathConstraint("wb_dma_infact_4par_seq_fields_cov_bin_scheme$__unbinned_filter");
        m_t2_channel_ac.setSpecificationComplete();
        m_path_coverages.push_back(m_t2_channel_ac);


        
        m_t3_channel_ac = new("t3.channel", {inst_name, "t3_channel_ac"}, eng);
        m_t3_channel_ac.addPathStopNode("t3.channel");
        m_t3_channel_ac.setGoalPathHitCount(1);
        m_t3_channel_ac.addBinScheme("wb_dma_infact_4par_seq_fields_cov_bin_scheme");
        m_t3_channel_ac.addPathConstraint("wb_dma_infact_4par_seq_fields_cov_bin_scheme$__unbinned_filter");
        m_t3_channel_ac.setSpecificationComplete();
        m_path_coverages.push_back(m_t3_channel_ac);


        
        m_t4_channel_ac = new("t4.channel", {inst_name, "t4_channel_ac"}, eng);
        m_t4_channel_ac.addPathStopNode("t4.channel");
        m_t4_channel_ac.setGoalPathHitCount(1);
        m_t4_channel_ac.addBinScheme("wb_dma_infact_4par_seq_fields_cov_bin_scheme");
        m_t4_channel_ac.addPathConstraint("wb_dma_infact_4par_seq_fields_cov_bin_scheme$__unbinned_filter");
        m_t4_channel_ac.setSpecificationComplete();
        m_path_coverages.push_back(m_t4_channel_ac);



	endfunction

	
 

       

	virtual function void delete();
		for (int i=0; i<m_path_coverages.size(); i++) begin
			m_path_coverages[i].delete();
		end
	endfunction 

	
 

	virtual function void getPathCoverageList(ref PathCoverage pc_list[$]);
		pc_list = m_path_coverages;
	endfunction

	
 

        

	virtual function void setPathCoverageCallback(PathCoverageCallback cb);
		for (int i=0; i<m_path_coverages.size(); i++) begin
			m_path_coverages[i].setCallback(cb);
		end
	endfunction

	
 

          
 

	virtual function void attach(TestEngine eng);
		for (int i=0; i<m_path_coverages.size(); i++) begin
			m_path_coverages[i].attach(eng);
		end
	endfunction 

	
 

          
 

	virtual function void detach(TestEngine eng);
		for (int i=0; i<m_path_coverages.size(); i++) begin
			m_path_coverages[i].detach(eng);
		end
	endfunction 

	
 

          
   

	virtual function bit allCoverageGoalsHaveBeenMet();
		bit ret = 1;
		for (int i=0; i<m_path_coverages.size(); i++) begin
			if (!m_path_coverages[i].allCoverageGoalsHaveBeenMet()) begin
				ret = 0;
				break;
			end
		end
		
		return ret;
	endfunction

	
 

          
      

	virtual function void setPriority(int base);
        m_t1_channel_ac.setPriority(base);
        m_t2_channel_ac.setPriority(base);
        m_t3_channel_ac.setPriority(base);
        m_t4_channel_ac.setPriority(base);

	endfunction

	
 

	virtual function string getCoverageReport();
		string report;
		int numTotal, numCov;
		bit allCount, allDone;
		
		report = $psprintf("%s\n%s\n%s\n",
			"---------------------------------------------------------------------",
			$psprintf("- wb_dma_infact_4par_seq_fields_cov Coverage Report: \"%s\"", m_inst_name),
			"---------------------------------------------------------------------");

		for (int i=0; i<m_path_coverages.size(); i++) begin
			allCount = m_path_coverages[i].currentResults(numTotal, numCov);
			allDone = m_path_coverages[i].allCoverageGoalsHaveBeenMet();
			report = {report, 
			$psprintf("    Path Coverage %0s: %0d/%0d%0s paths covered%0s\n",
				m_path_coverages[i].name(), numCov, numTotal, (allCount)?"":"+",
				(allDone)?" [COMPLETE]":"")};
		end

		return report;
	endfunction


endclass

 
`line 204 "wb_dma_infact_4par_seq_fields_cov.svh" 0
  


`line 206 "wb_dma_infact_4par_seq.svh" 0

  
`line 1 "wb_dma_infact_4par_seq_ll_single_cov.svh" 0

`line 1 "wb_dma_infact_4par_seq_ll_single_cov.svh" 0

 

        

       

  
`line 8 "wb_dma_infact_4par_seq_ll_single_cov.svh" 0

  
`line 9 "wb_dma_infact_4par_seq_ll_single_cov.svh" 0




class wb_dma_infact_4par_seq_ll_single_cov;

	
	
	
    PathCoverage                m_ll_size;




	
	PathCoverage						m_path_coverages[$];
	
	string								m_inst_name;

	

	
 

    

	function new(TestEngine eng, string inst_name="", bit instantiate_fc=1);
		string basename = inst_name;
		if (inst_name != "") begin
			inst_name = {inst_name, "."};
			m_inst_name = inst_name;
		end else begin
			m_inst_name = "";
		end
		
		if (instantiate_fc) begin

		end
        
        m_ll_size = new("do_4par", {inst_name, "ll_size"}, eng);
        m_ll_size.addPathStopNode("do_4par");
        m_ll_size.addBinScheme("ll_desc_sizes");
        m_ll_size.addPathConstraint("ll_desc_sizes$__unbinned_filter");
        m_ll_size.addBinScheme("dont_care$__t1.channel");
        m_ll_size.addBinScheme("dont_care$__t1.chk_sz");
        m_ll_size.addBinScheme("dont_care$__t1.dst_sel");
        m_ll_size.addBinScheme("dont_care$__t1.inc_dst");
        m_ll_size.addBinScheme("dont_care$__t1.inc_src");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[0].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[0].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[0].inc_src");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[0].src_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[0].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[10].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[10].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[10].inc_src");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[10].src_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[10].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[11].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[11].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[11].inc_src");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[11].src_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[11].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[12].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[12].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[12].inc_src");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[12].src_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[12].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[13].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[13].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[13].inc_src");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[13].src_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[13].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[14].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[14].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[14].inc_src");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[14].src_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[14].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[15].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[15].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[15].inc_src");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[15].src_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[15].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[1].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[1].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[1].inc_src");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[1].src_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[1].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[2].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[2].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[2].inc_src");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[2].src_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[2].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[3].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[3].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[3].inc_src");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[3].src_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[3].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[4].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[4].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[4].inc_src");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[4].src_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[4].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[5].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[5].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[5].inc_src");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[5].src_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[5].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[6].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[6].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[6].inc_src");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[6].src_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[6].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[7].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[7].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[7].inc_src");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[7].src_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[7].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[8].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[8].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[8].inc_src");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[8].src_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[8].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[9].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[9].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[9].inc_src");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[9].src_sel");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc[9].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc_tot_sz.sum");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc_tot_sz[0]");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc_tot_sz[10]");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc_tot_sz[11]");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc_tot_sz[12]");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc_tot_sz[13]");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc_tot_sz[14]");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc_tot_sz[15]");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc_tot_sz[1]");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc_tot_sz[2]");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc_tot_sz[3]");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc_tot_sz[4]");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc_tot_sz[5]");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc_tot_sz[6]");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc_tot_sz[7]");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc_tot_sz[8]");
        m_ll_size.addBinScheme("dont_care$__t1.ll_desc_tot_sz[9]");
        m_ll_size.addBinScheme("dont_care$__t1.mode");
        m_ll_size.addBinScheme("dont_care$__t1.src_sel");
        m_ll_size.addBinScheme("dont_care$__t1.tot_sz");
        m_ll_size.addBinScheme("dont_care$__t1.transfer_sz");
        m_ll_size.addBinScheme("dont_care$__t2.channel");
        m_ll_size.addBinScheme("dont_care$__t2.chk_sz");
        m_ll_size.addBinScheme("dont_care$__t2.dst_sel");
        m_ll_size.addBinScheme("dont_care$__t2.inc_dst");
        m_ll_size.addBinScheme("dont_care$__t2.inc_src");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[0].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[0].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[0].inc_src");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[0].src_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[0].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[10].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[10].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[10].inc_src");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[10].src_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[10].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[11].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[11].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[11].inc_src");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[11].src_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[11].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[12].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[12].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[12].inc_src");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[12].src_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[12].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[13].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[13].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[13].inc_src");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[13].src_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[13].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[14].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[14].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[14].inc_src");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[14].src_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[14].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[15].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[15].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[15].inc_src");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[15].src_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[15].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[1].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[1].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[1].inc_src");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[1].src_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[1].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[2].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[2].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[2].inc_src");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[2].src_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[2].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[3].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[3].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[3].inc_src");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[3].src_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[3].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[4].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[4].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[4].inc_src");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[4].src_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[4].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[5].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[5].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[5].inc_src");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[5].src_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[5].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[6].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[6].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[6].inc_src");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[6].src_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[6].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[7].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[7].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[7].inc_src");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[7].src_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[7].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[8].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[8].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[8].inc_src");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[8].src_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[8].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[9].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[9].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[9].inc_src");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[9].src_sel");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc[9].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc_tot_sz.sum");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc_tot_sz[0]");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc_tot_sz[10]");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc_tot_sz[11]");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc_tot_sz[12]");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc_tot_sz[13]");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc_tot_sz[14]");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc_tot_sz[15]");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc_tot_sz[1]");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc_tot_sz[2]");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc_tot_sz[3]");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc_tot_sz[4]");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc_tot_sz[5]");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc_tot_sz[6]");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc_tot_sz[7]");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc_tot_sz[8]");
        m_ll_size.addBinScheme("dont_care$__t2.ll_desc_tot_sz[9]");
        m_ll_size.addBinScheme("dont_care$__t2.mode");
        m_ll_size.addBinScheme("dont_care$__t2.src_sel");
        m_ll_size.addBinScheme("dont_care$__t2.tot_sz");
        m_ll_size.addBinScheme("dont_care$__t2.transfer_sz");
        m_ll_size.addBinScheme("dont_care$__t3.channel");
        m_ll_size.addBinScheme("dont_care$__t3.chk_sz");
        m_ll_size.addBinScheme("dont_care$__t3.dst_sel");
        m_ll_size.addBinScheme("dont_care$__t3.inc_dst");
        m_ll_size.addBinScheme("dont_care$__t3.inc_src");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[0].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[0].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[0].inc_src");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[0].src_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[0].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[10].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[10].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[10].inc_src");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[10].src_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[10].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[11].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[11].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[11].inc_src");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[11].src_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[11].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[12].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[12].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[12].inc_src");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[12].src_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[12].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[13].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[13].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[13].inc_src");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[13].src_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[13].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[14].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[14].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[14].inc_src");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[14].src_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[14].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[15].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[15].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[15].inc_src");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[15].src_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[15].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[1].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[1].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[1].inc_src");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[1].src_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[1].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[2].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[2].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[2].inc_src");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[2].src_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[2].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[3].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[3].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[3].inc_src");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[3].src_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[3].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[4].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[4].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[4].inc_src");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[4].src_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[4].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[5].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[5].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[5].inc_src");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[5].src_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[5].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[6].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[6].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[6].inc_src");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[6].src_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[6].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[7].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[7].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[7].inc_src");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[7].src_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[7].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[8].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[8].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[8].inc_src");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[8].src_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[8].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[9].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[9].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[9].inc_src");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[9].src_sel");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc[9].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc_tot_sz.sum");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc_tot_sz[0]");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc_tot_sz[10]");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc_tot_sz[11]");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc_tot_sz[12]");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc_tot_sz[13]");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc_tot_sz[14]");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc_tot_sz[15]");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc_tot_sz[1]");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc_tot_sz[2]");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc_tot_sz[3]");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc_tot_sz[4]");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc_tot_sz[5]");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc_tot_sz[6]");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc_tot_sz[7]");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc_tot_sz[8]");
        m_ll_size.addBinScheme("dont_care$__t3.ll_desc_tot_sz[9]");
        m_ll_size.addBinScheme("dont_care$__t3.mode");
        m_ll_size.addBinScheme("dont_care$__t3.src_sel");
        m_ll_size.addBinScheme("dont_care$__t3.tot_sz");
        m_ll_size.addBinScheme("dont_care$__t3.transfer_sz");
        m_ll_size.addBinScheme("dont_care$__t4.channel");
        m_ll_size.addBinScheme("dont_care$__t4.chk_sz");
        m_ll_size.addBinScheme("dont_care$__t4.dst_sel");
        m_ll_size.addBinScheme("dont_care$__t4.inc_dst");
        m_ll_size.addBinScheme("dont_care$__t4.inc_src");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[0].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[0].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[0].inc_src");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[0].src_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[0].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[10].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[10].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[10].inc_src");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[10].src_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[10].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[11].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[11].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[11].inc_src");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[11].src_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[11].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[12].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[12].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[12].inc_src");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[12].src_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[12].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[13].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[13].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[13].inc_src");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[13].src_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[13].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[14].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[14].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[14].inc_src");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[14].src_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[14].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[15].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[15].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[15].inc_src");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[15].src_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[15].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[1].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[1].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[1].inc_src");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[1].src_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[1].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[2].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[2].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[2].inc_src");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[2].src_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[2].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[3].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[3].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[3].inc_src");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[3].src_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[3].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[4].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[4].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[4].inc_src");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[4].src_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[4].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[5].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[5].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[5].inc_src");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[5].src_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[5].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[6].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[6].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[6].inc_src");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[6].src_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[6].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[7].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[7].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[7].inc_src");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[7].src_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[7].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[8].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[8].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[8].inc_src");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[8].src_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[8].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[9].dst_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[9].inc_dst");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[9].inc_src");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[9].src_sel");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc[9].tot_sz");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc_tot_sz.sum");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc_tot_sz[0]");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc_tot_sz[10]");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc_tot_sz[11]");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc_tot_sz[12]");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc_tot_sz[13]");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc_tot_sz[14]");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc_tot_sz[15]");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc_tot_sz[1]");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc_tot_sz[2]");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc_tot_sz[3]");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc_tot_sz[4]");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc_tot_sz[5]");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc_tot_sz[6]");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc_tot_sz[7]");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc_tot_sz[8]");
        m_ll_size.addBinScheme("dont_care$__t4.ll_desc_tot_sz[9]");
        m_ll_size.addBinScheme("dont_care$__t4.mode");
        m_ll_size.addBinScheme("dont_care$__t4.src_sel");
        m_ll_size.addBinScheme("dont_care$__t4.tot_sz");
        m_ll_size.addBinScheme("dont_care$__t4.transfer_sz");
        m_ll_size.setSpecificationComplete();
        m_path_coverages.push_back(m_ll_size);



	endfunction

	
 

       

	virtual function void delete();
		for (int i=0; i<m_path_coverages.size(); i++) begin
			m_path_coverages[i].delete();
		end
	endfunction 

	
 

	virtual function void getPathCoverageList(ref PathCoverage pc_list[$]);
		pc_list = m_path_coverages;
	endfunction

	
 

        

	virtual function void setPathCoverageCallback(PathCoverageCallback cb);
		for (int i=0; i<m_path_coverages.size(); i++) begin
			m_path_coverages[i].setCallback(cb);
		end
	endfunction

	
 

          
 

	virtual function void attach(TestEngine eng);
		for (int i=0; i<m_path_coverages.size(); i++) begin
			m_path_coverages[i].attach(eng);
		end
	endfunction 

	
 

          
 

	virtual function void detach(TestEngine eng);
		for (int i=0; i<m_path_coverages.size(); i++) begin
			m_path_coverages[i].detach(eng);
		end
	endfunction 

	
 

          
   

	virtual function bit allCoverageGoalsHaveBeenMet();
		bit ret = 1;
		for (int i=0; i<m_path_coverages.size(); i++) begin
			if (!m_path_coverages[i].allCoverageGoalsHaveBeenMet()) begin
				ret = 0;
				break;
			end
		end
		
		return ret;
	endfunction

	
 

          
      

	virtual function void setPriority(int base);
        m_ll_size.setPriority(base);

	endfunction

	
 

	virtual function string getCoverageReport();
		string report;
		int numTotal, numCov;
		bit allCount, allDone;
		
		report = $psprintf("%s\n%s\n%s\n",
			"---------------------------------------------------------------------",
			$psprintf("- wb_dma_infact_4par_seq_ll_single_cov Coverage Report: \"%s\"", m_inst_name),
			"---------------------------------------------------------------------");

		for (int i=0; i<m_path_coverages.size(); i++) begin
			allCount = m_path_coverages[i].currentResults(numTotal, numCov);
			allDone = m_path_coverages[i].allCoverageGoalsHaveBeenMet();
			report = {report, 
			$psprintf("    Path Coverage %0s: %0d/%0d%0s paths covered%0s\n",
				m_path_coverages[i].name(), numCov, numTotal, (allCount)?"":"+",
				(allDone)?" [COMPLETE]":"")};
		end

		return report;
	endfunction


endclass

 
`line 593 "wb_dma_infact_4par_seq_ll_single_cov.svh" 0
  


`line 595 "wb_dma_infact_4par_seq.svh" 0




  
`line 1 "wb_dma_infact_4par_seq_callback_closures.svh" 0

`line 1 "wb_dma_infact_4par_seq_callback_closures.svh" 0

 

        

       




class wb_dma_infact_4par_seq_pc_closure #(type T=int) extends PathCoverageCallback;
	T			m_target;
	
	function new(T target);
		m_target = target;
	endfunction
	
	virtual function void trigger(PathCoverage pc, CoverageCallbackReason reason);
		m_target.pathCoverageCallback(pc, reason);
	endfunction
	
endclass


`line 24 "wb_dma_infact_4par_seq.svh" 0


  
 
 
 
          
   










typedef wb_dma_multixfer_vseq wb_dma_infact_4par_seq_base_t;



typedef class wb_dma_infact_4par_seq_cb;




class wb_dma_infact_4par_seq extends wb_dma_infact_4par_seq_base_t;

    
	
    typedef wb_dma_infact_4par_seq wb_dma_infact_4par_seq_t;

    
     (

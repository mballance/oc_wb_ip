/****************************************************************************
 * wb_periph_subsys_w.sv
 ****************************************************************************/

/**
 * Module: wb_periph_subsys_w
 * 
 * Wire-based interface to the wb_periph_subsys module
 * 
 */
module wb_periph_subsys_w;


endmodule



/****************************************************************************
 * wb_simple_pic_dev_pkg.sv
 ****************************************************************************/
`include "uvm_macros.svh"
`include "uvmdev_macros.svh"

/**
 * Package: wb_simple_pic_dev_pkg
 * 
 * TODO: Add package documentation
 */
package wb_simple_pic_dev_pkg;
	import uvm_pkg::*;
	import uvmdev_pkg::*;
	import wb_simple_pic_reg_pkg::*;
	
	`include "wb_simple_pic_dev.svh"


endpackage




`include "uvm_macros.svh"

package wb_periph_subsys_env_pkg;
	import uvm_pkg::*;
	import wb_master_agent_pkg::*;
	import uart_serial_agent_pkg::*;
	import event_agent_pkg::*;

	`include "wb_periph_subsys_env.svh"
	
endpackage

/****************************************************************************
 * wb_uart_sequences_pkg.sv
 ****************************************************************************/

`include "uvm_macros.svh"

/**
 * Package: wb_uart_sequences_pkg
 * 
 * TODO: Add package documentation
 */
package wb_uart_sequences_pkg;
	import uvm_pkg::*;

	`include "wb_uart_vseq_base.svh"

endpackage



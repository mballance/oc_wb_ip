/****************************************************************************
 * wb_uart_dev_pkg.sv
 ****************************************************************************/
`include "uvm_macros.svh"
`include "uvmdev_macros.svh"

/**
 * Package: wb_uart_dev_pkg
 * 
 * TODO: Add package documentation
 */
package wb_uart_dev_pkg;
	import uvm_pkg::*;
	import uvmdev_pkg::*;
	import wb_uart_regs_pkg::*;
	
	`include "wb_uart_dev.svh"


endpackage



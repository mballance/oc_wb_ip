
`include "uvm_macros.svh"

package wb_periph_subsys_env_pkg;
	import uvm_pkg::*;

	`include "wb_periph_subsys_env.svh"
	
endpackage

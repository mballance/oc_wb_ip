/****************************************************************************
 * wb_periph_subsys_seqs_pkg.sv
 ****************************************************************************/
`include "uvm_macros.svh"

/**
 * Package: wb_periph_subsys_seqs_pkg
 * 
 * TODO: Add package documentation
 */
package wb_periph_subsys_seqs_pkg;
	import uvm_pkg::*;
	
	`include "wb_periph_subsys_vseq.svh"


endpackage



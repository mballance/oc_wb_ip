
`include "uvm_macros.svh"

package wb_uart_env_pkg;
	import uvm_pkg::*;

	`include "wb_uart_env.svh"
	
endpackage
